`define CROSSBAR_INST(n) \
    axi_crossbar_``n`` axi_crossbar_inst ( \
        .aclk(aclk), \
        .aresetn(aresetn), \
        .s_axi_awid(s_axi_awid), \
        .s_axi_awaddr(s_axi_awaddr), \
        .s_axi_awlen(s_axi_awlen), \
        .s_axi_awsize(s_axi_awsize), \
        .s_axi_awburst(s_axi_awburst), \
        .s_axi_awlock(s_axi_awlock), \
        .s_axi_awcache(s_axi_awcache), \
        .s_axi_awprot(s_axi_awprot), \
        .s_axi_awqos(s_axi_awqos), \
        .s_axi_awvalid(s_axi_awvalid), \
        .s_axi_awready(s_axi_awready), \
        .s_axi_wdata(s_axi_wdata), \
        .s_axi_wstrb(s_axi_wstrb), \
        .s_axi_wlast(s_axi_wlast), \
        .s_axi_wvalid(s_axi_wvalid), \
        .s_axi_wready(s_axi_wready), \
        .s_axi_bid(s_axi_bid), \
        .s_axi_bresp(s_axi_bresp), \
        .s_axi_bvalid(s_axi_bvalid), \
        .s_axi_bready(s_axi_bready), \
        .s_axi_arid(s_axi_arid), \
        .s_axi_araddr(s_axi_araddr), \
        .s_axi_arlen(s_axi_arlen), \
        .s_axi_arsize(s_axi_arsize), \
        .s_axi_arburst(s_axi_arburst), \
        .s_axi_arlock(s_axi_arlock), \
        .s_axi_arcache(s_axi_arcache), \
        .s_axi_arprot(s_axi_arprot), \
        .s_axi_arqos(s_axi_arqos), \
        .s_axi_arvalid(s_axi_arvalid), \
        .s_axi_arready(s_axi_arready), \
        .s_axi_rid(s_axi_rid), \
        .s_axi_rdata(s_axi_rdata), \
        .s_axi_rresp(s_axi_rresp), \
        .s_axi_rlast(s_axi_rlast), \
        .s_axi_rvalid(s_axi_rvalid), \
        .s_axi_rready(s_axi_rready), \
        .m_axi_awid(m_axi_awid), \
        .m_axi_awaddr(m_axi_awaddr), \
        .m_axi_awlen(m_axi_awlen), \
        .m_axi_awsize(m_axi_awsize), \
        .m_axi_awburst(m_axi_awburst), \
        .m_axi_awlock(m_axi_awlock), \
        .m_axi_awcache(m_axi_awcache), \
        .m_axi_awprot(m_axi_awprot), \
        .m_axi_awregion(m_axi_awregion), \
        .m_axi_awqos(m_axi_awqos), \
        .m_axi_awvalid(m_axi_awvalid), \
        .m_axi_awready(m_axi_awready), \
        .m_axi_wdata(m_axi_wdata), \
        .m_axi_wstrb(m_axi_wstrb), \
        .m_axi_wlast(m_axi_wlast), \
        .m_axi_wvalid(m_axi_wvalid), \
        .m_axi_wready(m_axi_wready), \
        .m_axi_bid(m_axi_bid), \
        .m_axi_bresp(m_axi_bresp), \
        .m_axi_bvalid(m_axi_bvalid), \
        .m_axi_bready(m_axi_bready), \
        .m_axi_arid(m_axi_arid), \
        .m_axi_araddr(m_axi_araddr), \
        .m_axi_arlen(m_axi_arlen), \
        .m_axi_arsize(m_axi_arsize), \
        .m_axi_arburst(m_axi_arburst), \
        .m_axi_arlock(m_axi_arlock), \
        .m_axi_arcache(m_axi_arcache), \
        .m_axi_arprot(m_axi_arprot), \
        .m_axi_arregion(m_axi_arregion), \
        .m_axi_arqos(m_axi_arqos), \
        .m_axi_arvalid(m_axi_arvalid), \
        .m_axi_arready(m_axi_arready), \
        .m_axi_rid(m_axi_rid), \
        .m_axi_rdata(m_axi_rdata), \
        .m_axi_rresp(m_axi_rresp), \
        .m_axi_rlast(m_axi_rlast), \
        .m_axi_rvalid(m_axi_rvalid), \
        .m_axi_rready(m_axi_rready) \
    );

`define AXI_PORT_LIST(n) \
    input wire [ID_WIDTH-1 : 0] s_axi_``n``_awid, \
    input wire [(32*1)-1 : 0] s_axi_``n``_awaddr, \
    input wire [(8*1)-1 : 0] s_axi_``n``_awlen, \
    input wire [(3*1)-1 : 0] s_axi_``n``_awsize, \
    input wire [(2*1)-1 : 0] s_axi_``n``_awburst, \
    input wire [1-1 : 0] s_axi_``n``_awlock, \
    input wire [(4*1)-1 : 0] s_axi_``n``_awcache, \
    input wire [(3*1)-1 : 0] s_axi_``n``_awprot, \
    input wire [(4*1)-1 : 0] s_axi_``n``_awqos, \
    input wire [1-1 : 0] s_axi_``n``_awvalid, \
    output wire [1-1 : 0] s_axi_``n``_awready, \
    input wire [(64*1)-1 : 0] s_axi_``n``_wdata, \
    input wire [(8*1)-1 : 0] s_axi_``n``_wstrb, \
    input wire [1-1 : 0] s_axi_``n``_wlast, \
    input wire [1-1 : 0] s_axi_``n``_wvalid, \
    output wire [1-1 : 0] s_axi_``n``_wready, \
    output wire [ID_WIDTH-1 : 0] s_axi_``n``_bid, \
    output wire [(2*1)-1 : 0] s_axi_``n``_bresp, \
    output wire [1-1 : 0] s_axi_``n``_bvalid, \
    input wire [1-1 : 0] s_axi_``n``_bready, \
    input wire [ID_WIDTH-1 : 0] s_axi_``n``_arid, \
    input wire [(32*1)-1 : 0] s_axi_``n``_araddr, \
    input wire [(8*1)-1 : 0] s_axi_``n``_arlen, \
    input wire [(3*1)-1 : 0] s_axi_``n``_arsize, \
    input wire [(2*1)-1 : 0] s_axi_``n``_arburst, \
    input wire [1-1 : 0] s_axi_``n``_arlock, \
    input wire [(4*1)-1 : 0] s_axi_``n``_arcache, \
    input wire [(3*1)-1 : 0] s_axi_``n``_arprot, \
    input wire [(4*1)-1 : 0] s_axi_``n``_arqos, \
    input wire [1-1 : 0] s_axi_``n``_arvalid, \
    output wire [1-1 : 0] s_axi_``n``_arready, \
    output wire [ID_WIDTH-1 : 0] s_axi_``n``_rid, \
    output wire [(64*1)-1 : 0] s_axi_``n``_rdata, \
    output wire [(2*1)-1 : 0] s_axi_``n``_rresp, \
    output wire [1-1 : 0] s_axi_``n``_rlast, \
    output wire [1-1 : 0] s_axi_``n``_rvalid, \
    input wire [1-1 : 0] s_axi_``n``_rready

module memory #(
    parameter KERNELS = 16,
    parameter ID_WIDTH = KERNELS == 1 ? 1 : $clog2(KERNELS)
)(
    input wire aclk,
    input wire aresetn,

    `AXI_PORT_LIST(0),
    `AXI_PORT_LIST(1),
    `AXI_PORT_LIST(2),
    `AXI_PORT_LIST(3),
    `AXI_PORT_LIST(4),
    `AXI_PORT_LIST(5),
    `AXI_PORT_LIST(6),
    `AXI_PORT_LIST(7),
    `AXI_PORT_LIST(8),
    `AXI_PORT_LIST(9),
    `AXI_PORT_LIST(10),
    `AXI_PORT_LIST(11),
    `AXI_PORT_LIST(12),
    `AXI_PORT_LIST(13),
    `AXI_PORT_LIST(14),
    `AXI_PORT_LIST(15),    

    output wire [ID_WIDTH-1 : 0] m_axi_awid,
    output wire [31 : 0] m_axi_awaddr,
    output wire [7 : 0] m_axi_awlen,
    output wire [2 : 0] m_axi_awsize,
    output wire [1 : 0] m_axi_awburst,
    output wire [0 : 0] m_axi_awlock,
    output wire [3 : 0] m_axi_awcache,
    output wire [2 : 0] m_axi_awprot,
    output wire [3 : 0] m_axi_awregion,
    output wire [3 : 0] m_axi_awqos,
    output wire [0 : 0] m_axi_awvalid,
    input wire [0 : 0] m_axi_awready,
    output wire [63 : 0] m_axi_wdata,
    output wire [7 : 0] m_axi_wstrb,
    output wire [0 : 0] m_axi_wlast,
    output wire [0 : 0] m_axi_wvalid,
    input wire [0 : 0] m_axi_wready,
    input wire [ID_WIDTH-1 : 0] m_axi_bid,
    input wire [1 : 0] m_axi_bresp,
    input wire [0 : 0] m_axi_bvalid,
    output wire [0 : 0] m_axi_bready,
    output wire [ID_WIDTH-1 : 0] m_axi_arid,
    output wire [31 : 0] m_axi_araddr,
    output wire [7 : 0] m_axi_arlen,
    output wire [2 : 0] m_axi_arsize,
    output wire [1 : 0] m_axi_arburst,
    output wire [0 : 0] m_axi_arlock,
    output wire [3 : 0] m_axi_arcache,
    output wire [2 : 0] m_axi_arprot,
    output wire [3 : 0] m_axi_arregion,
    output wire [3 : 0] m_axi_arqos,
    output wire [0 : 0] m_axi_arvalid,
    input wire [0 : 0] m_axi_arready,
    input wire [ID_WIDTH-1 : 0] m_axi_rid,
    input wire [63 : 0] m_axi_rdata,
    input wire [1 : 0] m_axi_rresp,
    input wire [0 : 0] m_axi_rlast,
    input wire [0 : 0] m_axi_rvalid,
    output wire [0 : 0] m_axi_rready
);

wire [(ID_WIDTH*KERNELS)-1 : 0] s_axi_awid;
wire [(32*KERNELS)-1 : 0] s_axi_awaddr;
wire [(8*KERNELS)-1 : 0] s_axi_awlen;
wire [(3*KERNELS)-1 : 0] s_axi_awsize;
wire [(2*KERNELS)-1 : 0] s_axi_awburst;
wire [KERNELS-1 : 0] s_axi_awlock;
wire [(4*KERNELS)-1 : 0] s_axi_awcache;
wire [(3*KERNELS)-1 : 0] s_axi_awprot;
wire [(4*KERNELS)-1 : 0] s_axi_awqos;
wire [KERNELS-1 : 0] s_axi_awvalid;
wire [KERNELS-1 : 0] s_axi_awready;
wire [(64*KERNELS)-1 : 0] s_axi_wdata;
wire [(8*KERNELS)-1 : 0] s_axi_wstrb;
wire [KERNELS-1 : 0] s_axi_wlast;
wire [KERNELS-1 : 0] s_axi_wvalid;
wire [KERNELS-1 : 0] s_axi_wready;
wire [(ID_WIDTH*KERNELS)-1 : 0] s_axi_bid;
wire [(2*KERNELS)-1 : 0] s_axi_bresp;
wire [KERNELS-1 : 0] s_axi_bvalid;
wire [KERNELS-1 : 0] s_axi_bready;
wire [(ID_WIDTH*KERNELS)-1 : 0] s_axi_arid;
wire [(32*KERNELS)-1 : 0] s_axi_araddr;
wire [(8*KERNELS)-1 : 0] s_axi_arlen;
wire [(3*KERNELS)-1 : 0] s_axi_arsize;
wire [(2*KERNELS)-1 : 0] s_axi_arburst;
wire [KERNELS-1 : 0] s_axi_arlock;
wire [(4*KERNELS)-1 : 0] s_axi_arcache;
wire [(3*KERNELS)-1 : 0] s_axi_arprot;
wire [(4*KERNELS)-1 : 0] s_axi_arqos;
wire [KERNELS-1 : 0] s_axi_arvalid;
wire [KERNELS-1 : 0] s_axi_arready;
wire [(ID_WIDTH*KERNELS)-1 : 0] s_axi_rid;
wire [(64*KERNELS)-1 : 0] s_axi_rdata;
wire [(2*KERNELS)-1 : 0] s_axi_rresp;
wire [KERNELS-1 : 0] s_axi_rlast;
wire [KERNELS-1 : 0] s_axi_rvalid;
wire [KERNELS-1 : 0] s_axi_rready;

generate
    case(KERNELS)
        1: begin
            assign s_axi_awid = s_axi_0_awid;
            assign s_axi_awaddr = s_axi_0_awaddr;
            assign s_axi_awlen = s_axi_0_awlen;
            assign s_axi_awsize = s_axi_0_awsize;
            assign s_axi_awburst = s_axi_0_awburst;
            assign s_axi_awlock = s_axi_0_awlock;
            assign s_axi_awcache = s_axi_0_awcache;
            assign s_axi_awprot = s_axi_0_awprot;
            assign s_axi_awqos = s_axi_0_awqos;
            assign s_axi_awvalid = s_axi_0_awvalid;
            assign s_axi_0_awready = s_axi_awready;
            assign s_axi_wdata = s_axi_0_wdata;
            assign s_axi_wstrb = s_axi_0_wstrb;
            assign s_axi_wlast = s_axi_0_wlast;
            assign s_axi_wvalid = s_axi_0_wvalid;
            assign s_axi_0_wready = s_axi_wready;
            assign s_axi_0_bid = s_axi_bid;
            assign s_axi_0_bresp = s_axi_bresp;
            assign s_axi_0_bvalid = s_axi_bvalid;
            assign s_axi_bready = s_axi_0_bready;
            assign s_axi_arid = s_axi_0_arid;
            assign s_axi_araddr = s_axi_0_araddr;
            assign s_axi_arlen = s_axi_0_arlen;
            assign s_axi_arsize = s_axi_0_arsize;
            assign s_axi_arburst = s_axi_0_arburst;
            assign s_axi_arlock = s_axi_0_arlock;
            assign s_axi_arcache = s_axi_0_arcache;
            assign s_axi_arprot = s_axi_0_arprot;
            assign s_axi_arqos = s_axi_0_arqos;
            assign s_axi_arvalid = s_axi_0_arvalid;
            assign s_axi_0_arready = s_axi_arready;
            assign s_axi_0_rid = s_axi_rid;
            assign s_axi_0_rdata = s_axi_rdata;
            assign s_axi_0_rresp = s_axi_rresp;
            assign s_axi_0_rlast = s_axi_rlast;
            assign s_axi_0_rvalid = s_axi_rvalid;
            assign s_axi_rready = s_axi_0_rready;
        end
        2: begin
            assign s_axi_awid = {s_axi_1_awid,s_axi_0_awid};
            assign s_axi_awaddr = {s_axi_1_awaddr,s_axi_0_awaddr};
            assign s_axi_awlen = {s_axi_1_awlen,s_axi_0_awlen};
            assign s_axi_awsize = {s_axi_1_awsize,s_axi_0_awsize};
            assign s_axi_awburst = {s_axi_1_awburst,s_axi_0_awburst};
            assign s_axi_awlock = {s_axi_1_awlock,s_axi_0_awlock};
            assign s_axi_awcache = {s_axi_1_awcache,s_axi_0_awcache};
            assign s_axi_awprot = {s_axi_1_awprot,s_axi_0_awprot};
            assign s_axi_awqos = {s_axi_1_awqos,s_axi_0_awqos};
            assign s_axi_awvalid = {s_axi_1_awvalid,s_axi_0_awvalid};
            assign {s_axi_1_awready,s_axi_0_awready} = s_axi_awready;
            assign s_axi_wdata = {s_axi_1_wdata,s_axi_0_wdata};
            assign s_axi_wstrb = {s_axi_1_wstrb,s_axi_0_wstrb};
            assign s_axi_wlast = {s_axi_1_wlast,s_axi_0_wlast};
            assign s_axi_wvalid = {s_axi_1_wvalid,s_axi_0_wvalid};
            assign {s_axi_1_wready,s_axi_0_wready} = s_axi_wready;
            assign {s_axi_1_bid,s_axi_0_bid} = s_axi_bid;
            assign {s_axi_1_bresp,s_axi_0_bresp} = s_axi_bresp;
            assign {s_axi_1_bvalid,s_axi_0_bvalid} = s_axi_bvalid;
            assign s_axi_bready = {s_axi_1_bready,s_axi_0_bready};
            assign s_axi_arid = {s_axi_1_arid,s_axi_0_arid};
            assign s_axi_araddr = {s_axi_1_araddr,s_axi_0_araddr};
            assign s_axi_arlen = {s_axi_1_arlen,s_axi_0_arlen};
            assign s_axi_arsize = {s_axi_1_arsize,s_axi_0_arsize};
            assign s_axi_arburst = {s_axi_1_arburst,s_axi_0_arburst};
            assign s_axi_arlock = {s_axi_1_arlock,s_axi_0_arlock};
            assign s_axi_arcache = {s_axi_1_arcache,s_axi_0_arcache};
            assign s_axi_arprot = {s_axi_1_arprot,s_axi_0_arprot};
            assign s_axi_arqos = {s_axi_1_arqos,s_axi_0_arqos};
            assign s_axi_arvalid = {s_axi_1_arvalid,s_axi_0_arvalid};
            assign {s_axi_1_arready,s_axi_0_arready} = s_axi_arready;
            assign {s_axi_1_rid,s_axi_0_rid} = s_axi_rid;
            assign {s_axi_1_rdata,s_axi_0_rdata} = s_axi_rdata;
            assign {s_axi_1_rresp,s_axi_0_rresp} = s_axi_rresp;
            assign {s_axi_1_rlast,s_axi_0_rlast} = s_axi_rlast;
            assign {s_axi_1_rvalid,s_axi_0_rvalid} = s_axi_rvalid;
            assign s_axi_rready = {s_axi_1_rready,s_axi_0_rready};
        end
        3: begin
            assign s_axi_awid = {s_axi_2_awid,s_axi_1_awid,s_axi_0_awid};
            assign s_axi_awaddr = {s_axi_2_awaddr,s_axi_1_awaddr,s_axi_0_awaddr};
            assign s_axi_awlen = {s_axi_2_awlen,s_axi_1_awlen,s_axi_0_awlen};
            assign s_axi_awsize = {s_axi_2_awsize,s_axi_1_awsize,s_axi_0_awsize};
            assign s_axi_awburst = {s_axi_2_awburst,s_axi_1_awburst,s_axi_0_awburst};
            assign s_axi_awlock = {s_axi_2_awlock,s_axi_1_awlock,s_axi_0_awlock};
            assign s_axi_awcache = {s_axi_2_awcache,s_axi_1_awcache,s_axi_0_awcache};
            assign s_axi_awprot = {s_axi_2_awprot,s_axi_1_awprot,s_axi_0_awprot};
            assign s_axi_awqos = {s_axi_2_awqos,s_axi_1_awqos,s_axi_0_awqos};
            assign s_axi_awvalid = {s_axi_2_awvalid,s_axi_1_awvalid,s_axi_0_awvalid};
            assign {s_axi_2_awready,s_axi_1_awready,s_axi_0_awready} = s_axi_awready;
            assign s_axi_wdata = {s_axi_2_wdata,s_axi_1_wdata,s_axi_0_wdata};
            assign s_axi_wstrb = {s_axi_2_wstrb,s_axi_1_wstrb,s_axi_0_wstrb};
            assign s_axi_wlast = {s_axi_2_wlast,s_axi_1_wlast,s_axi_0_wlast};
            assign s_axi_wvalid = {s_axi_2_wvalid,s_axi_1_wvalid,s_axi_0_wvalid};
            assign {s_axi_2_wready,s_axi_1_wready,s_axi_0_wready} = s_axi_wready;
            assign {s_axi_2_bid,s_axi_1_bid,s_axi_0_bid} = s_axi_bid;
            assign {s_axi_2_bresp,s_axi_1_bresp,s_axi_0_bresp} = s_axi_bresp;
            assign {s_axi_2_bvalid,s_axi_1_bvalid,s_axi_0_bvalid} = s_axi_bvalid;
            assign s_axi_bready = {s_axi_2_bready,s_axi_1_bready,s_axi_0_bready};
            assign s_axi_arid = {s_axi_2_arid,s_axi_1_arid,s_axi_0_arid};
            assign s_axi_araddr = {s_axi_2_araddr,s_axi_1_araddr,s_axi_0_araddr};
            assign s_axi_arlen = {s_axi_2_arlen,s_axi_1_arlen,s_axi_0_arlen};
            assign s_axi_arsize = {s_axi_2_arsize,s_axi_1_arsize,s_axi_0_arsize};
            assign s_axi_arburst = {s_axi_2_arburst,s_axi_1_arburst,s_axi_0_arburst};
            assign s_axi_arlock = {s_axi_2_arlock,s_axi_1_arlock,s_axi_0_arlock};
            assign s_axi_arcache = {s_axi_2_arcache,s_axi_1_arcache,s_axi_0_arcache};
            assign s_axi_arprot = {s_axi_2_arprot,s_axi_1_arprot,s_axi_0_arprot};
            assign s_axi_arqos = {s_axi_2_arqos,s_axi_1_arqos,s_axi_0_arqos};
            assign s_axi_arvalid = {s_axi_2_arvalid,s_axi_1_arvalid,s_axi_0_arvalid};
            assign {s_axi_2_arready,s_axi_1_arready,s_axi_0_arready} = s_axi_arready;
            assign {s_axi_2_rid,s_axi_1_rid,s_axi_0_rid} = s_axi_rid;
            assign {s_axi_2_rdata,s_axi_1_rdata,s_axi_0_rdata} = s_axi_rdata;
            assign {s_axi_2_rresp,s_axi_1_rresp,s_axi_0_rresp} = s_axi_rresp;
            assign {s_axi_2_rlast,s_axi_1_rlast,s_axi_0_rlast} = s_axi_rlast;
            assign {s_axi_2_rvalid,s_axi_1_rvalid,s_axi_0_rvalid} = s_axi_rvalid;
            assign s_axi_rready = {s_axi_2_rready,s_axi_1_rready,s_axi_0_rready};
        end
        4: begin
            assign s_axi_awid = {s_axi_3_awid,s_axi_2_awid,s_axi_1_awid,s_axi_0_awid};
            assign s_axi_awaddr = {s_axi_3_awaddr,s_axi_2_awaddr,s_axi_1_awaddr,s_axi_0_awaddr};
            assign s_axi_awlen = {s_axi_3_awlen,s_axi_2_awlen,s_axi_1_awlen,s_axi_0_awlen};
            assign s_axi_awsize = {s_axi_3_awsize,s_axi_2_awsize,s_axi_1_awsize,s_axi_0_awsize};
            assign s_axi_awburst = {s_axi_3_awburst,s_axi_2_awburst,s_axi_1_awburst,s_axi_0_awburst};
            assign s_axi_awlock = {s_axi_3_awlock,s_axi_2_awlock,s_axi_1_awlock,s_axi_0_awlock};
            assign s_axi_awcache = {s_axi_3_awcache,s_axi_2_awcache,s_axi_1_awcache,s_axi_0_awcache};
            assign s_axi_awprot = {s_axi_3_awprot,s_axi_2_awprot,s_axi_1_awprot,s_axi_0_awprot};
            assign s_axi_awqos = {s_axi_3_awqos,s_axi_2_awqos,s_axi_1_awqos,s_axi_0_awqos};
            assign s_axi_awvalid = {s_axi_3_awvalid,s_axi_2_awvalid,s_axi_1_awvalid,s_axi_0_awvalid};
            assign {s_axi_3_awready,s_axi_2_awready,s_axi_1_awready,s_axi_0_awready} = s_axi_awready;
            assign s_axi_wdata = {s_axi_3_wdata,s_axi_2_wdata,s_axi_1_wdata,s_axi_0_wdata};
            assign s_axi_wstrb = {s_axi_3_wstrb,s_axi_2_wstrb,s_axi_1_wstrb,s_axi_0_wstrb};
            assign s_axi_wlast = {s_axi_3_wlast,s_axi_2_wlast,s_axi_1_wlast,s_axi_0_wlast};
            assign s_axi_wvalid = {s_axi_3_wvalid,s_axi_2_wvalid,s_axi_1_wvalid,s_axi_0_wvalid};
            assign {s_axi_3_wready,s_axi_2_wready,s_axi_1_wready,s_axi_0_wready} = s_axi_wready;
            assign {s_axi_3_bid,s_axi_2_bid,s_axi_1_bid,s_axi_0_bid} = s_axi_bid;
            assign {s_axi_3_bresp,s_axi_2_bresp,s_axi_1_bresp,s_axi_0_bresp} = s_axi_bresp;
            assign {s_axi_3_bvalid,s_axi_2_bvalid,s_axi_1_bvalid,s_axi_0_bvalid} = s_axi_bvalid;
            assign s_axi_bready = {s_axi_3_bready,s_axi_2_bready,s_axi_1_bready,s_axi_0_bready};
            assign s_axi_arid = {s_axi_3_arid,s_axi_2_arid,s_axi_1_arid,s_axi_0_arid};
            assign s_axi_araddr = {s_axi_3_araddr,s_axi_2_araddr,s_axi_1_araddr,s_axi_0_araddr};
            assign s_axi_arlen = {s_axi_3_arlen,s_axi_2_arlen,s_axi_1_arlen,s_axi_0_arlen};
            assign s_axi_arsize = {s_axi_3_arsize,s_axi_2_arsize,s_axi_1_arsize,s_axi_0_arsize};
            assign s_axi_arburst = {s_axi_3_arburst,s_axi_2_arburst,s_axi_1_arburst,s_axi_0_arburst};
            assign s_axi_arlock = {s_axi_3_arlock,s_axi_2_arlock,s_axi_1_arlock,s_axi_0_arlock};
            assign s_axi_arcache = {s_axi_3_arcache,s_axi_2_arcache,s_axi_1_arcache,s_axi_0_arcache};
            assign s_axi_arprot = {s_axi_3_arprot,s_axi_2_arprot,s_axi_1_arprot,s_axi_0_arprot};
            assign s_axi_arqos = {s_axi_3_arqos,s_axi_2_arqos,s_axi_1_arqos,s_axi_0_arqos};
            assign s_axi_arvalid = {s_axi_3_arvalid,s_axi_2_arvalid,s_axi_1_arvalid,s_axi_0_arvalid};
            assign {s_axi_3_arready,s_axi_2_arready,s_axi_1_arready,s_axi_0_arready} = s_axi_arready;
            assign {s_axi_3_rid,s_axi_2_rid,s_axi_1_rid,s_axi_0_rid} = s_axi_rid;
            assign {s_axi_3_rdata,s_axi_2_rdata,s_axi_1_rdata,s_axi_0_rdata} = s_axi_rdata;
            assign {s_axi_3_rresp,s_axi_2_rresp,s_axi_1_rresp,s_axi_0_rresp} = s_axi_rresp;
            assign {s_axi_3_rlast,s_axi_2_rlast,s_axi_1_rlast,s_axi_0_rlast} = s_axi_rlast;
            assign {s_axi_3_rvalid,s_axi_2_rvalid,s_axi_1_rvalid,s_axi_0_rvalid} = s_axi_rvalid;
            assign s_axi_rready = {s_axi_3_rready,s_axi_2_rready,s_axi_1_rready,s_axi_0_rready};
        end
        5: begin
            assign s_axi_awid = {s_axi_4_awid,s_axi_3_awid,s_axi_2_awid,s_axi_1_awid,s_axi_0_awid};
            assign s_axi_awaddr = {s_axi_4_awaddr,s_axi_3_awaddr,s_axi_2_awaddr,s_axi_1_awaddr,s_axi_0_awaddr};
            assign s_axi_awlen = {s_axi_4_awlen,s_axi_3_awlen,s_axi_2_awlen,s_axi_1_awlen,s_axi_0_awlen};
            assign s_axi_awsize = {s_axi_4_awsize,s_axi_3_awsize,s_axi_2_awsize,s_axi_1_awsize,s_axi_0_awsize};
            assign s_axi_awburst = {s_axi_4_awburst,s_axi_3_awburst,s_axi_2_awburst,s_axi_1_awburst,s_axi_0_awburst};
            assign s_axi_awlock = {s_axi_4_awlock,s_axi_3_awlock,s_axi_2_awlock,s_axi_1_awlock,s_axi_0_awlock};
            assign s_axi_awcache = {s_axi_4_awcache,s_axi_3_awcache,s_axi_2_awcache,s_axi_1_awcache,s_axi_0_awcache};
            assign s_axi_awprot = {s_axi_4_awprot,s_axi_3_awprot,s_axi_2_awprot,s_axi_1_awprot,s_axi_0_awprot};
            assign s_axi_awqos = {s_axi_4_awqos,s_axi_3_awqos,s_axi_2_awqos,s_axi_1_awqos,s_axi_0_awqos};
            assign s_axi_awvalid = {s_axi_4_awvalid,s_axi_3_awvalid,s_axi_2_awvalid,s_axi_1_awvalid,s_axi_0_awvalid};
            assign {s_axi_4_awready,s_axi_3_awready,s_axi_2_awready,s_axi_1_awready,s_axi_0_awready} = s_axi_awready;
            assign s_axi_wdata = {s_axi_4_wdata,s_axi_3_wdata,s_axi_2_wdata,s_axi_1_wdata,s_axi_0_wdata};
            assign s_axi_wstrb = {s_axi_4_wstrb,s_axi_3_wstrb,s_axi_2_wstrb,s_axi_1_wstrb,s_axi_0_wstrb};
            assign s_axi_wlast = {s_axi_4_wlast,s_axi_3_wlast,s_axi_2_wlast,s_axi_1_wlast,s_axi_0_wlast};
            assign s_axi_wvalid = {s_axi_4_wvalid,s_axi_3_wvalid,s_axi_2_wvalid,s_axi_1_wvalid,s_axi_0_wvalid};
            assign {s_axi_4_wready,s_axi_3_wready,s_axi_2_wready,s_axi_1_wready,s_axi_0_wready} = s_axi_wready;
            assign {s_axi_4_bid,s_axi_3_bid,s_axi_2_bid,s_axi_1_bid,s_axi_0_bid} = s_axi_bid;
            assign {s_axi_4_bresp,s_axi_3_bresp,s_axi_2_bresp,s_axi_1_bresp,s_axi_0_bresp} = s_axi_bresp;
            assign {s_axi_4_bvalid,s_axi_3_bvalid,s_axi_2_bvalid,s_axi_1_bvalid,s_axi_0_bvalid} = s_axi_bvalid;
            assign s_axi_bready = {s_axi_4_bready,s_axi_3_bready,s_axi_2_bready,s_axi_1_bready,s_axi_0_bready};
            assign s_axi_arid = {s_axi_4_arid,s_axi_3_arid,s_axi_2_arid,s_axi_1_arid,s_axi_0_arid};
            assign s_axi_araddr = {s_axi_4_araddr,s_axi_3_araddr,s_axi_2_araddr,s_axi_1_araddr,s_axi_0_araddr};
            assign s_axi_arlen = {s_axi_4_arlen,s_axi_3_arlen,s_axi_2_arlen,s_axi_1_arlen,s_axi_0_arlen};
            assign s_axi_arsize = {s_axi_4_arsize,s_axi_3_arsize,s_axi_2_arsize,s_axi_1_arsize,s_axi_0_arsize};
            assign s_axi_arburst = {s_axi_4_arburst,s_axi_3_arburst,s_axi_2_arburst,s_axi_1_arburst,s_axi_0_arburst};
            assign s_axi_arlock = {s_axi_4_arlock,s_axi_3_arlock,s_axi_2_arlock,s_axi_1_arlock,s_axi_0_arlock};
            assign s_axi_arcache = {s_axi_4_arcache,s_axi_3_arcache,s_axi_2_arcache,s_axi_1_arcache,s_axi_0_arcache};
            assign s_axi_arprot = {s_axi_4_arprot,s_axi_3_arprot,s_axi_2_arprot,s_axi_1_arprot,s_axi_0_arprot};
            assign s_axi_arqos = {s_axi_4_arqos,s_axi_3_arqos,s_axi_2_arqos,s_axi_1_arqos,s_axi_0_arqos};
            assign s_axi_arvalid = {s_axi_4_arvalid,s_axi_3_arvalid,s_axi_2_arvalid,s_axi_1_arvalid,s_axi_0_arvalid};
            assign {s_axi_4_arready,s_axi_3_arready,s_axi_2_arready,s_axi_1_arready,s_axi_0_arready} = s_axi_arready;
            assign {s_axi_4_rid,s_axi_3_rid,s_axi_2_rid,s_axi_1_rid,s_axi_0_rid} = s_axi_rid;
            assign {s_axi_4_rdata,s_axi_3_rdata,s_axi_2_rdata,s_axi_1_rdata,s_axi_0_rdata} = s_axi_rdata;
            assign {s_axi_4_rresp,s_axi_3_rresp,s_axi_2_rresp,s_axi_1_rresp,s_axi_0_rresp} = s_axi_rresp;
            assign {s_axi_4_rlast,s_axi_3_rlast,s_axi_2_rlast,s_axi_1_rlast,s_axi_0_rlast} = s_axi_rlast;
            assign {s_axi_4_rvalid,s_axi_3_rvalid,s_axi_2_rvalid,s_axi_1_rvalid,s_axi_0_rvalid} = s_axi_rvalid;
            assign s_axi_rready = {s_axi_4_rready,s_axi_3_rready,s_axi_2_rready,s_axi_1_rready,s_axi_0_rready};
        end
        6: begin
            assign s_axi_awid = {s_axi_5_awid,s_axi_4_awid,s_axi_3_awid,s_axi_2_awid,s_axi_1_awid,s_axi_0_awid};
            assign s_axi_awaddr = {s_axi_5_awaddr,s_axi_4_awaddr,s_axi_3_awaddr,s_axi_2_awaddr,s_axi_1_awaddr,s_axi_0_awaddr};
            assign s_axi_awlen = {s_axi_5_awlen,s_axi_4_awlen,s_axi_3_awlen,s_axi_2_awlen,s_axi_1_awlen,s_axi_0_awlen};
            assign s_axi_awsize = {s_axi_5_awsize,s_axi_4_awsize,s_axi_3_awsize,s_axi_2_awsize,s_axi_1_awsize,s_axi_0_awsize};
            assign s_axi_awburst = {s_axi_5_awburst,s_axi_4_awburst,s_axi_3_awburst,s_axi_2_awburst,s_axi_1_awburst,s_axi_0_awburst};
            assign s_axi_awlock = {s_axi_5_awlock,s_axi_4_awlock,s_axi_3_awlock,s_axi_2_awlock,s_axi_1_awlock,s_axi_0_awlock};
            assign s_axi_awcache = {s_axi_5_awcache,s_axi_4_awcache,s_axi_3_awcache,s_axi_2_awcache,s_axi_1_awcache,s_axi_0_awcache};
            assign s_axi_awprot = {s_axi_5_awprot,s_axi_4_awprot,s_axi_3_awprot,s_axi_2_awprot,s_axi_1_awprot,s_axi_0_awprot};
            assign s_axi_awqos = {s_axi_5_awqos,s_axi_4_awqos,s_axi_3_awqos,s_axi_2_awqos,s_axi_1_awqos,s_axi_0_awqos};
            assign s_axi_awvalid = {s_axi_5_awvalid,s_axi_4_awvalid,s_axi_3_awvalid,s_axi_2_awvalid,s_axi_1_awvalid,s_axi_0_awvalid};
            assign {s_axi_5_awready,s_axi_4_awready,s_axi_3_awready,s_axi_2_awready,s_axi_1_awready,s_axi_0_awready} = s_axi_awready;
            assign s_axi_wdata = {s_axi_5_wdata,s_axi_4_wdata,s_axi_3_wdata,s_axi_2_wdata,s_axi_1_wdata,s_axi_0_wdata};
            assign s_axi_wstrb = {s_axi_5_wstrb,s_axi_4_wstrb,s_axi_3_wstrb,s_axi_2_wstrb,s_axi_1_wstrb,s_axi_0_wstrb};
            assign s_axi_wlast = {s_axi_5_wlast,s_axi_4_wlast,s_axi_3_wlast,s_axi_2_wlast,s_axi_1_wlast,s_axi_0_wlast};
            assign s_axi_wvalid = {s_axi_5_wvalid,s_axi_4_wvalid,s_axi_3_wvalid,s_axi_2_wvalid,s_axi_1_wvalid,s_axi_0_wvalid};
            assign {s_axi_5_wready,s_axi_4_wready,s_axi_3_wready,s_axi_2_wready,s_axi_1_wready,s_axi_0_wready} = s_axi_wready;
            assign {s_axi_5_bid,s_axi_4_bid,s_axi_3_bid,s_axi_2_bid,s_axi_1_bid,s_axi_0_bid} = s_axi_bid;
            assign {s_axi_5_bresp,s_axi_4_bresp,s_axi_3_bresp,s_axi_2_bresp,s_axi_1_bresp,s_axi_0_bresp} = s_axi_bresp;
            assign {s_axi_5_bvalid,s_axi_4_bvalid,s_axi_3_bvalid,s_axi_2_bvalid,s_axi_1_bvalid,s_axi_0_bvalid} = s_axi_bvalid;
            assign s_axi_bready = {s_axi_5_bready,s_axi_4_bready,s_axi_3_bready,s_axi_2_bready,s_axi_1_bready,s_axi_0_bready};
            assign s_axi_arid = {s_axi_5_arid,s_axi_4_arid,s_axi_3_arid,s_axi_2_arid,s_axi_1_arid,s_axi_0_arid};
            assign s_axi_araddr = {s_axi_5_araddr,s_axi_4_araddr,s_axi_3_araddr,s_axi_2_araddr,s_axi_1_araddr,s_axi_0_araddr};
            assign s_axi_arlen = {s_axi_5_arlen,s_axi_4_arlen,s_axi_3_arlen,s_axi_2_arlen,s_axi_1_arlen,s_axi_0_arlen};
            assign s_axi_arsize = {s_axi_5_arsize,s_axi_4_arsize,s_axi_3_arsize,s_axi_2_arsize,s_axi_1_arsize,s_axi_0_arsize};
            assign s_axi_arburst = {s_axi_5_arburst,s_axi_4_arburst,s_axi_3_arburst,s_axi_2_arburst,s_axi_1_arburst,s_axi_0_arburst};
            assign s_axi_arlock = {s_axi_5_arlock,s_axi_4_arlock,s_axi_3_arlock,s_axi_2_arlock,s_axi_1_arlock,s_axi_0_arlock};
            assign s_axi_arcache = {s_axi_5_arcache,s_axi_4_arcache,s_axi_3_arcache,s_axi_2_arcache,s_axi_1_arcache,s_axi_0_arcache};
            assign s_axi_arprot = {s_axi_5_arprot,s_axi_4_arprot,s_axi_3_arprot,s_axi_2_arprot,s_axi_1_arprot,s_axi_0_arprot};
            assign s_axi_arqos = {s_axi_5_arqos,s_axi_4_arqos,s_axi_3_arqos,s_axi_2_arqos,s_axi_1_arqos,s_axi_0_arqos};
            assign s_axi_arvalid = {s_axi_5_arvalid,s_axi_4_arvalid,s_axi_3_arvalid,s_axi_2_arvalid,s_axi_1_arvalid,s_axi_0_arvalid};
            assign {s_axi_5_arready,s_axi_4_arready,s_axi_3_arready,s_axi_2_arready,s_axi_1_arready,s_axi_0_arready} = s_axi_arready;
            assign {s_axi_5_rid,s_axi_4_rid,s_axi_3_rid,s_axi_2_rid,s_axi_1_rid,s_axi_0_rid} = s_axi_rid;
            assign {s_axi_5_rdata,s_axi_4_rdata,s_axi_3_rdata,s_axi_2_rdata,s_axi_1_rdata,s_axi_0_rdata} = s_axi_rdata;
            assign {s_axi_5_rresp,s_axi_4_rresp,s_axi_3_rresp,s_axi_2_rresp,s_axi_1_rresp,s_axi_0_rresp} = s_axi_rresp;
            assign {s_axi_5_rlast,s_axi_4_rlast,s_axi_3_rlast,s_axi_2_rlast,s_axi_1_rlast,s_axi_0_rlast} = s_axi_rlast;
            assign {s_axi_5_rvalid,s_axi_4_rvalid,s_axi_3_rvalid,s_axi_2_rvalid,s_axi_1_rvalid,s_axi_0_rvalid} = s_axi_rvalid;
            assign s_axi_rready = {s_axi_5_rready,s_axi_4_rready,s_axi_3_rready,s_axi_2_rready,s_axi_1_rready,s_axi_0_rready};
        end
        7: begin
            assign s_axi_awid = {s_axi_6_awid,s_axi_5_awid,s_axi_4_awid,s_axi_3_awid,s_axi_2_awid,s_axi_1_awid,s_axi_0_awid};
            assign s_axi_awaddr = {s_axi_6_awaddr,s_axi_5_awaddr,s_axi_4_awaddr,s_axi_3_awaddr,s_axi_2_awaddr,s_axi_1_awaddr,s_axi_0_awaddr};
            assign s_axi_awlen = {s_axi_6_awlen,s_axi_5_awlen,s_axi_4_awlen,s_axi_3_awlen,s_axi_2_awlen,s_axi_1_awlen,s_axi_0_awlen};
            assign s_axi_awsize = {s_axi_6_awsize,s_axi_5_awsize,s_axi_4_awsize,s_axi_3_awsize,s_axi_2_awsize,s_axi_1_awsize,s_axi_0_awsize};
            assign s_axi_awburst = {s_axi_6_awburst,s_axi_5_awburst,s_axi_4_awburst,s_axi_3_awburst,s_axi_2_awburst,s_axi_1_awburst,s_axi_0_awburst};
            assign s_axi_awlock = {s_axi_6_awlock,s_axi_5_awlock,s_axi_4_awlock,s_axi_3_awlock,s_axi_2_awlock,s_axi_1_awlock,s_axi_0_awlock};
            assign s_axi_awcache = {s_axi_6_awcache,s_axi_5_awcache,s_axi_4_awcache,s_axi_3_awcache,s_axi_2_awcache,s_axi_1_awcache,s_axi_0_awcache};
            assign s_axi_awprot = {s_axi_6_awprot,s_axi_5_awprot,s_axi_4_awprot,s_axi_3_awprot,s_axi_2_awprot,s_axi_1_awprot,s_axi_0_awprot};
            assign s_axi_awqos = {s_axi_6_awqos,s_axi_5_awqos,s_axi_4_awqos,s_axi_3_awqos,s_axi_2_awqos,s_axi_1_awqos,s_axi_0_awqos};
            assign s_axi_awvalid = {s_axi_6_awvalid,s_axi_5_awvalid,s_axi_4_awvalid,s_axi_3_awvalid,s_axi_2_awvalid,s_axi_1_awvalid,s_axi_0_awvalid};
            assign {s_axi_6_awready,s_axi_5_awready,s_axi_4_awready,s_axi_3_awready,s_axi_2_awready,s_axi_1_awready,s_axi_0_awready} = s_axi_awready;
            assign s_axi_wdata = {s_axi_6_wdata,s_axi_5_wdata,s_axi_4_wdata,s_axi_3_wdata,s_axi_2_wdata,s_axi_1_wdata,s_axi_0_wdata};
            assign s_axi_wstrb = {s_axi_6_wstrb,s_axi_5_wstrb,s_axi_4_wstrb,s_axi_3_wstrb,s_axi_2_wstrb,s_axi_1_wstrb,s_axi_0_wstrb};
            assign s_axi_wlast = {s_axi_6_wlast,s_axi_5_wlast,s_axi_4_wlast,s_axi_3_wlast,s_axi_2_wlast,s_axi_1_wlast,s_axi_0_wlast};
            assign s_axi_wvalid = {s_axi_6_wvalid,s_axi_5_wvalid,s_axi_4_wvalid,s_axi_3_wvalid,s_axi_2_wvalid,s_axi_1_wvalid,s_axi_0_wvalid};
            assign {s_axi_6_wready,s_axi_5_wready,s_axi_4_wready,s_axi_3_wready,s_axi_2_wready,s_axi_1_wready,s_axi_0_wready} = s_axi_wready;
            assign {s_axi_6_bid,s_axi_5_bid,s_axi_4_bid,s_axi_3_bid,s_axi_2_bid,s_axi_1_bid,s_axi_0_bid} = s_axi_bid;
            assign {s_axi_6_bresp,s_axi_5_bresp,s_axi_4_bresp,s_axi_3_bresp,s_axi_2_bresp,s_axi_1_bresp,s_axi_0_bresp} = s_axi_bresp;
            assign {s_axi_6_bvalid,s_axi_5_bvalid,s_axi_4_bvalid,s_axi_3_bvalid,s_axi_2_bvalid,s_axi_1_bvalid,s_axi_0_bvalid} = s_axi_bvalid;
            assign s_axi_bready = {s_axi_6_bready,s_axi_5_bready,s_axi_4_bready,s_axi_3_bready,s_axi_2_bready,s_axi_1_bready,s_axi_0_bready};
            assign s_axi_arid = {s_axi_6_arid,s_axi_5_arid,s_axi_4_arid,s_axi_3_arid,s_axi_2_arid,s_axi_1_arid,s_axi_0_arid};
            assign s_axi_araddr = {s_axi_6_araddr,s_axi_5_araddr,s_axi_4_araddr,s_axi_3_araddr,s_axi_2_araddr,s_axi_1_araddr,s_axi_0_araddr};
            assign s_axi_arlen = {s_axi_6_arlen,s_axi_5_arlen,s_axi_4_arlen,s_axi_3_arlen,s_axi_2_arlen,s_axi_1_arlen,s_axi_0_arlen};
            assign s_axi_arsize = {s_axi_6_arsize,s_axi_5_arsize,s_axi_4_arsize,s_axi_3_arsize,s_axi_2_arsize,s_axi_1_arsize,s_axi_0_arsize};
            assign s_axi_arburst = {s_axi_6_arburst,s_axi_5_arburst,s_axi_4_arburst,s_axi_3_arburst,s_axi_2_arburst,s_axi_1_arburst,s_axi_0_arburst};
            assign s_axi_arlock = {s_axi_6_arlock,s_axi_5_arlock,s_axi_4_arlock,s_axi_3_arlock,s_axi_2_arlock,s_axi_1_arlock,s_axi_0_arlock};
            assign s_axi_arcache = {s_axi_6_arcache,s_axi_5_arcache,s_axi_4_arcache,s_axi_3_arcache,s_axi_2_arcache,s_axi_1_arcache,s_axi_0_arcache};
            assign s_axi_arprot = {s_axi_6_arprot,s_axi_5_arprot,s_axi_4_arprot,s_axi_3_arprot,s_axi_2_arprot,s_axi_1_arprot,s_axi_0_arprot};
            assign s_axi_arqos = {s_axi_6_arqos,s_axi_5_arqos,s_axi_4_arqos,s_axi_3_arqos,s_axi_2_arqos,s_axi_1_arqos,s_axi_0_arqos};
            assign s_axi_arvalid = {s_axi_6_arvalid,s_axi_5_arvalid,s_axi_4_arvalid,s_axi_3_arvalid,s_axi_2_arvalid,s_axi_1_arvalid,s_axi_0_arvalid};
            assign {s_axi_6_arready,s_axi_5_arready,s_axi_4_arready,s_axi_3_arready,s_axi_2_arready,s_axi_1_arready,s_axi_0_arready} = s_axi_arready;
            assign {s_axi_6_rid,s_axi_5_rid,s_axi_4_rid,s_axi_3_rid,s_axi_2_rid,s_axi_1_rid,s_axi_0_rid} = s_axi_rid;
            assign {s_axi_6_rdata,s_axi_5_rdata,s_axi_4_rdata,s_axi_3_rdata,s_axi_2_rdata,s_axi_1_rdata,s_axi_0_rdata} = s_axi_rdata;
            assign {s_axi_6_rresp,s_axi_5_rresp,s_axi_4_rresp,s_axi_3_rresp,s_axi_2_rresp,s_axi_1_rresp,s_axi_0_rresp} = s_axi_rresp;
            assign {s_axi_6_rlast,s_axi_5_rlast,s_axi_4_rlast,s_axi_3_rlast,s_axi_2_rlast,s_axi_1_rlast,s_axi_0_rlast} = s_axi_rlast;
            assign {s_axi_6_rvalid,s_axi_5_rvalid,s_axi_4_rvalid,s_axi_3_rvalid,s_axi_2_rvalid,s_axi_1_rvalid,s_axi_0_rvalid} = s_axi_rvalid;
            assign s_axi_rready = {s_axi_6_rready,s_axi_5_rready,s_axi_4_rready,s_axi_3_rready,s_axi_2_rready,s_axi_1_rready,s_axi_0_rready};
        end
        8: begin
            assign s_axi_awid = {s_axi_7_awid,s_axi_6_awid,s_axi_5_awid,s_axi_4_awid,s_axi_3_awid,s_axi_2_awid,s_axi_1_awid,s_axi_0_awid};
            assign s_axi_awaddr = {s_axi_7_awaddr,s_axi_6_awaddr,s_axi_5_awaddr,s_axi_4_awaddr,s_axi_3_awaddr,s_axi_2_awaddr,s_axi_1_awaddr,s_axi_0_awaddr};
            assign s_axi_awlen = {s_axi_7_awlen,s_axi_6_awlen,s_axi_5_awlen,s_axi_4_awlen,s_axi_3_awlen,s_axi_2_awlen,s_axi_1_awlen,s_axi_0_awlen};
            assign s_axi_awsize = {s_axi_7_awsize,s_axi_6_awsize,s_axi_5_awsize,s_axi_4_awsize,s_axi_3_awsize,s_axi_2_awsize,s_axi_1_awsize,s_axi_0_awsize};
            assign s_axi_awburst = {s_axi_7_awburst,s_axi_6_awburst,s_axi_5_awburst,s_axi_4_awburst,s_axi_3_awburst,s_axi_2_awburst,s_axi_1_awburst,s_axi_0_awburst};
            assign s_axi_awlock = {s_axi_7_awlock,s_axi_6_awlock,s_axi_5_awlock,s_axi_4_awlock,s_axi_3_awlock,s_axi_2_awlock,s_axi_1_awlock,s_axi_0_awlock};
            assign s_axi_awcache = {s_axi_7_awcache,s_axi_6_awcache,s_axi_5_awcache,s_axi_4_awcache,s_axi_3_awcache,s_axi_2_awcache,s_axi_1_awcache,s_axi_0_awcache};
            assign s_axi_awprot = {s_axi_7_awprot,s_axi_6_awprot,s_axi_5_awprot,s_axi_4_awprot,s_axi_3_awprot,s_axi_2_awprot,s_axi_1_awprot,s_axi_0_awprot};
            assign s_axi_awqos = {s_axi_7_awqos,s_axi_6_awqos,s_axi_5_awqos,s_axi_4_awqos,s_axi_3_awqos,s_axi_2_awqos,s_axi_1_awqos,s_axi_0_awqos};
            assign s_axi_awvalid = {s_axi_7_awvalid,s_axi_6_awvalid,s_axi_5_awvalid,s_axi_4_awvalid,s_axi_3_awvalid,s_axi_2_awvalid,s_axi_1_awvalid,s_axi_0_awvalid};
            assign {s_axi_7_awready,s_axi_6_awready,s_axi_5_awready,s_axi_4_awready,s_axi_3_awready,s_axi_2_awready,s_axi_1_awready,s_axi_0_awready} = s_axi_awready;
            assign s_axi_wdata = {s_axi_7_wdata,s_axi_6_wdata,s_axi_5_wdata,s_axi_4_wdata,s_axi_3_wdata,s_axi_2_wdata,s_axi_1_wdata,s_axi_0_wdata};
            assign s_axi_wstrb = {s_axi_7_wstrb,s_axi_6_wstrb,s_axi_5_wstrb,s_axi_4_wstrb,s_axi_3_wstrb,s_axi_2_wstrb,s_axi_1_wstrb,s_axi_0_wstrb};
            assign s_axi_wlast = {s_axi_7_wlast,s_axi_6_wlast,s_axi_5_wlast,s_axi_4_wlast,s_axi_3_wlast,s_axi_2_wlast,s_axi_1_wlast,s_axi_0_wlast};
            assign s_axi_wvalid = {s_axi_7_wvalid,s_axi_6_wvalid,s_axi_5_wvalid,s_axi_4_wvalid,s_axi_3_wvalid,s_axi_2_wvalid,s_axi_1_wvalid,s_axi_0_wvalid};
            assign {s_axi_7_wready,s_axi_6_wready,s_axi_5_wready,s_axi_4_wready,s_axi_3_wready,s_axi_2_wready,s_axi_1_wready,s_axi_0_wready} = s_axi_wready;
            assign {s_axi_7_bid,s_axi_6_bid,s_axi_5_bid,s_axi_4_bid,s_axi_3_bid,s_axi_2_bid,s_axi_1_bid,s_axi_0_bid} = s_axi_bid;
            assign {s_axi_7_bresp,s_axi_6_bresp,s_axi_5_bresp,s_axi_4_bresp,s_axi_3_bresp,s_axi_2_bresp,s_axi_1_bresp,s_axi_0_bresp} = s_axi_bresp;
            assign {s_axi_7_bvalid,s_axi_6_bvalid,s_axi_5_bvalid,s_axi_4_bvalid,s_axi_3_bvalid,s_axi_2_bvalid,s_axi_1_bvalid,s_axi_0_bvalid} = s_axi_bvalid;
            assign s_axi_bready = {s_axi_7_bready,s_axi_6_bready,s_axi_5_bready,s_axi_4_bready,s_axi_3_bready,s_axi_2_bready,s_axi_1_bready,s_axi_0_bready};
            assign s_axi_arid = {s_axi_7_arid,s_axi_6_arid,s_axi_5_arid,s_axi_4_arid,s_axi_3_arid,s_axi_2_arid,s_axi_1_arid,s_axi_0_arid};
            assign s_axi_araddr = {s_axi_7_araddr,s_axi_6_araddr,s_axi_5_araddr,s_axi_4_araddr,s_axi_3_araddr,s_axi_2_araddr,s_axi_1_araddr,s_axi_0_araddr};
            assign s_axi_arlen = {s_axi_7_arlen,s_axi_6_arlen,s_axi_5_arlen,s_axi_4_arlen,s_axi_3_arlen,s_axi_2_arlen,s_axi_1_arlen,s_axi_0_arlen};
            assign s_axi_arsize = {s_axi_7_arsize,s_axi_6_arsize,s_axi_5_arsize,s_axi_4_arsize,s_axi_3_arsize,s_axi_2_arsize,s_axi_1_arsize,s_axi_0_arsize};
            assign s_axi_arburst = {s_axi_7_arburst,s_axi_6_arburst,s_axi_5_arburst,s_axi_4_arburst,s_axi_3_arburst,s_axi_2_arburst,s_axi_1_arburst,s_axi_0_arburst};
            assign s_axi_arlock = {s_axi_7_arlock,s_axi_6_arlock,s_axi_5_arlock,s_axi_4_arlock,s_axi_3_arlock,s_axi_2_arlock,s_axi_1_arlock,s_axi_0_arlock};
            assign s_axi_arcache = {s_axi_7_arcache,s_axi_6_arcache,s_axi_5_arcache,s_axi_4_arcache,s_axi_3_arcache,s_axi_2_arcache,s_axi_1_arcache,s_axi_0_arcache};
            assign s_axi_arprot = {s_axi_7_arprot,s_axi_6_arprot,s_axi_5_arprot,s_axi_4_arprot,s_axi_3_arprot,s_axi_2_arprot,s_axi_1_arprot,s_axi_0_arprot};
            assign s_axi_arqos = {s_axi_7_arqos,s_axi_6_arqos,s_axi_5_arqos,s_axi_4_arqos,s_axi_3_arqos,s_axi_2_arqos,s_axi_1_arqos,s_axi_0_arqos};
            assign s_axi_arvalid = {s_axi_7_arvalid,s_axi_6_arvalid,s_axi_5_arvalid,s_axi_4_arvalid,s_axi_3_arvalid,s_axi_2_arvalid,s_axi_1_arvalid,s_axi_0_arvalid};
            assign {s_axi_7_arready,s_axi_6_arready,s_axi_5_arready,s_axi_4_arready,s_axi_3_arready,s_axi_2_arready,s_axi_1_arready,s_axi_0_arready} = s_axi_arready;
            assign {s_axi_7_rid,s_axi_6_rid,s_axi_5_rid,s_axi_4_rid,s_axi_3_rid,s_axi_2_rid,s_axi_1_rid,s_axi_0_rid} = s_axi_rid;
            assign {s_axi_7_rdata,s_axi_6_rdata,s_axi_5_rdata,s_axi_4_rdata,s_axi_3_rdata,s_axi_2_rdata,s_axi_1_rdata,s_axi_0_rdata} = s_axi_rdata;
            assign {s_axi_7_rresp,s_axi_6_rresp,s_axi_5_rresp,s_axi_4_rresp,s_axi_3_rresp,s_axi_2_rresp,s_axi_1_rresp,s_axi_0_rresp} = s_axi_rresp;
            assign {s_axi_7_rlast,s_axi_6_rlast,s_axi_5_rlast,s_axi_4_rlast,s_axi_3_rlast,s_axi_2_rlast,s_axi_1_rlast,s_axi_0_rlast} = s_axi_rlast;
            assign {s_axi_7_rvalid,s_axi_6_rvalid,s_axi_5_rvalid,s_axi_4_rvalid,s_axi_3_rvalid,s_axi_2_rvalid,s_axi_1_rvalid,s_axi_0_rvalid} = s_axi_rvalid;
            assign s_axi_rready = {s_axi_7_rready,s_axi_6_rready,s_axi_5_rready,s_axi_4_rready,s_axi_3_rready,s_axi_2_rready,s_axi_1_rready,s_axi_0_rready};
        end
        9: begin
            assign s_axi_awid = {s_axi_8_awid,s_axi_7_awid,s_axi_6_awid,s_axi_5_awid,s_axi_4_awid,s_axi_3_awid,s_axi_2_awid,s_axi_1_awid,s_axi_0_awid};
            assign s_axi_awaddr = {s_axi_8_awaddr,s_axi_7_awaddr,s_axi_6_awaddr,s_axi_5_awaddr,s_axi_4_awaddr,s_axi_3_awaddr,s_axi_2_awaddr,s_axi_1_awaddr,s_axi_0_awaddr};
            assign s_axi_awlen = {s_axi_8_awlen,s_axi_7_awlen,s_axi_6_awlen,s_axi_5_awlen,s_axi_4_awlen,s_axi_3_awlen,s_axi_2_awlen,s_axi_1_awlen,s_axi_0_awlen};
            assign s_axi_awsize = {s_axi_8_awsize,s_axi_7_awsize,s_axi_6_awsize,s_axi_5_awsize,s_axi_4_awsize,s_axi_3_awsize,s_axi_2_awsize,s_axi_1_awsize,s_axi_0_awsize};
            assign s_axi_awburst = {s_axi_8_awburst,s_axi_7_awburst,s_axi_6_awburst,s_axi_5_awburst,s_axi_4_awburst,s_axi_3_awburst,s_axi_2_awburst,s_axi_1_awburst,s_axi_0_awburst};
            assign s_axi_awlock = {s_axi_8_awlock,s_axi_7_awlock,s_axi_6_awlock,s_axi_5_awlock,s_axi_4_awlock,s_axi_3_awlock,s_axi_2_awlock,s_axi_1_awlock,s_axi_0_awlock};
            assign s_axi_awcache = {s_axi_8_awcache,s_axi_7_awcache,s_axi_6_awcache,s_axi_5_awcache,s_axi_4_awcache,s_axi_3_awcache,s_axi_2_awcache,s_axi_1_awcache,s_axi_0_awcache};
            assign s_axi_awprot = {s_axi_8_awprot,s_axi_7_awprot,s_axi_6_awprot,s_axi_5_awprot,s_axi_4_awprot,s_axi_3_awprot,s_axi_2_awprot,s_axi_1_awprot,s_axi_0_awprot};
            assign s_axi_awqos = {s_axi_8_awqos,s_axi_7_awqos,s_axi_6_awqos,s_axi_5_awqos,s_axi_4_awqos,s_axi_3_awqos,s_axi_2_awqos,s_axi_1_awqos,s_axi_0_awqos};
            assign s_axi_awvalid = {s_axi_8_awvalid,s_axi_7_awvalid,s_axi_6_awvalid,s_axi_5_awvalid,s_axi_4_awvalid,s_axi_3_awvalid,s_axi_2_awvalid,s_axi_1_awvalid,s_axi_0_awvalid};
            assign {s_axi_8_awready,s_axi_7_awready,s_axi_6_awready,s_axi_5_awready,s_axi_4_awready,s_axi_3_awready,s_axi_2_awready,s_axi_1_awready,s_axi_0_awready} = s_axi_awready;
            assign s_axi_wdata = {s_axi_8_wdata,s_axi_7_wdata,s_axi_6_wdata,s_axi_5_wdata,s_axi_4_wdata,s_axi_3_wdata,s_axi_2_wdata,s_axi_1_wdata,s_axi_0_wdata};
            assign s_axi_wstrb = {s_axi_8_wstrb,s_axi_7_wstrb,s_axi_6_wstrb,s_axi_5_wstrb,s_axi_4_wstrb,s_axi_3_wstrb,s_axi_2_wstrb,s_axi_1_wstrb,s_axi_0_wstrb};
            assign s_axi_wlast = {s_axi_8_wlast,s_axi_7_wlast,s_axi_6_wlast,s_axi_5_wlast,s_axi_4_wlast,s_axi_3_wlast,s_axi_2_wlast,s_axi_1_wlast,s_axi_0_wlast};
            assign s_axi_wvalid = {s_axi_8_wvalid,s_axi_7_wvalid,s_axi_6_wvalid,s_axi_5_wvalid,s_axi_4_wvalid,s_axi_3_wvalid,s_axi_2_wvalid,s_axi_1_wvalid,s_axi_0_wvalid};
            assign {s_axi_8_wready,s_axi_7_wready,s_axi_6_wready,s_axi_5_wready,s_axi_4_wready,s_axi_3_wready,s_axi_2_wready,s_axi_1_wready,s_axi_0_wready} = s_axi_wready;
            assign {s_axi_8_bid,s_axi_7_bid,s_axi_6_bid,s_axi_5_bid,s_axi_4_bid,s_axi_3_bid,s_axi_2_bid,s_axi_1_bid,s_axi_0_bid} = s_axi_bid;
            assign {s_axi_8_bresp,s_axi_7_bresp,s_axi_6_bresp,s_axi_5_bresp,s_axi_4_bresp,s_axi_3_bresp,s_axi_2_bresp,s_axi_1_bresp,s_axi_0_bresp} = s_axi_bresp;
            assign {s_axi_8_bvalid,s_axi_7_bvalid,s_axi_6_bvalid,s_axi_5_bvalid,s_axi_4_bvalid,s_axi_3_bvalid,s_axi_2_bvalid,s_axi_1_bvalid,s_axi_0_bvalid} = s_axi_bvalid;
            assign s_axi_bready = {s_axi_8_bready,s_axi_7_bready,s_axi_6_bready,s_axi_5_bready,s_axi_4_bready,s_axi_3_bready,s_axi_2_bready,s_axi_1_bready,s_axi_0_bready};
            assign s_axi_arid = {s_axi_8_arid,s_axi_7_arid,s_axi_6_arid,s_axi_5_arid,s_axi_4_arid,s_axi_3_arid,s_axi_2_arid,s_axi_1_arid,s_axi_0_arid};
            assign s_axi_araddr = {s_axi_8_araddr,s_axi_7_araddr,s_axi_6_araddr,s_axi_5_araddr,s_axi_4_araddr,s_axi_3_araddr,s_axi_2_araddr,s_axi_1_araddr,s_axi_0_araddr};
            assign s_axi_arlen = {s_axi_8_arlen,s_axi_7_arlen,s_axi_6_arlen,s_axi_5_arlen,s_axi_4_arlen,s_axi_3_arlen,s_axi_2_arlen,s_axi_1_arlen,s_axi_0_arlen};
            assign s_axi_arsize = {s_axi_8_arsize,s_axi_7_arsize,s_axi_6_arsize,s_axi_5_arsize,s_axi_4_arsize,s_axi_3_arsize,s_axi_2_arsize,s_axi_1_arsize,s_axi_0_arsize};
            assign s_axi_arburst = {s_axi_8_arburst,s_axi_7_arburst,s_axi_6_arburst,s_axi_5_arburst,s_axi_4_arburst,s_axi_3_arburst,s_axi_2_arburst,s_axi_1_arburst,s_axi_0_arburst};
            assign s_axi_arlock = {s_axi_8_arlock,s_axi_7_arlock,s_axi_6_arlock,s_axi_5_arlock,s_axi_4_arlock,s_axi_3_arlock,s_axi_2_arlock,s_axi_1_arlock,s_axi_0_arlock};
            assign s_axi_arcache = {s_axi_8_arcache,s_axi_7_arcache,s_axi_6_arcache,s_axi_5_arcache,s_axi_4_arcache,s_axi_3_arcache,s_axi_2_arcache,s_axi_1_arcache,s_axi_0_arcache};
            assign s_axi_arprot = {s_axi_8_arprot,s_axi_7_arprot,s_axi_6_arprot,s_axi_5_arprot,s_axi_4_arprot,s_axi_3_arprot,s_axi_2_arprot,s_axi_1_arprot,s_axi_0_arprot};
            assign s_axi_arqos = {s_axi_8_arqos,s_axi_7_arqos,s_axi_6_arqos,s_axi_5_arqos,s_axi_4_arqos,s_axi_3_arqos,s_axi_2_arqos,s_axi_1_arqos,s_axi_0_arqos};
            assign s_axi_arvalid = {s_axi_8_arvalid,s_axi_7_arvalid,s_axi_6_arvalid,s_axi_5_arvalid,s_axi_4_arvalid,s_axi_3_arvalid,s_axi_2_arvalid,s_axi_1_arvalid,s_axi_0_arvalid};
            assign {s_axi_8_arready,s_axi_7_arready,s_axi_6_arready,s_axi_5_arready,s_axi_4_arready,s_axi_3_arready,s_axi_2_arready,s_axi_1_arready,s_axi_0_arready} = s_axi_arready;
            assign {s_axi_8_rid,s_axi_7_rid,s_axi_6_rid,s_axi_5_rid,s_axi_4_rid,s_axi_3_rid,s_axi_2_rid,s_axi_1_rid,s_axi_0_rid} = s_axi_rid;
            assign {s_axi_8_rdata,s_axi_7_rdata,s_axi_6_rdata,s_axi_5_rdata,s_axi_4_rdata,s_axi_3_rdata,s_axi_2_rdata,s_axi_1_rdata,s_axi_0_rdata} = s_axi_rdata;
            assign {s_axi_8_rresp,s_axi_7_rresp,s_axi_6_rresp,s_axi_5_rresp,s_axi_4_rresp,s_axi_3_rresp,s_axi_2_rresp,s_axi_1_rresp,s_axi_0_rresp} = s_axi_rresp;
            assign {s_axi_8_rlast,s_axi_7_rlast,s_axi_6_rlast,s_axi_5_rlast,s_axi_4_rlast,s_axi_3_rlast,s_axi_2_rlast,s_axi_1_rlast,s_axi_0_rlast} = s_axi_rlast;
            assign {s_axi_8_rvalid,s_axi_7_rvalid,s_axi_6_rvalid,s_axi_5_rvalid,s_axi_4_rvalid,s_axi_3_rvalid,s_axi_2_rvalid,s_axi_1_rvalid,s_axi_0_rvalid} = s_axi_rvalid;
            assign s_axi_rready = {s_axi_8_rready,s_axi_7_rready,s_axi_6_rready,s_axi_5_rready,s_axi_4_rready,s_axi_3_rready,s_axi_2_rready,s_axi_1_rready,s_axi_0_rready};
        end
        10: begin
            assign s_axi_awid = {s_axi_9_awid,s_axi_8_awid,s_axi_7_awid,s_axi_6_awid,s_axi_5_awid,s_axi_4_awid,s_axi_3_awid,s_axi_2_awid,s_axi_1_awid,s_axi_0_awid};
            assign s_axi_awaddr = {s_axi_9_awaddr,s_axi_8_awaddr,s_axi_7_awaddr,s_axi_6_awaddr,s_axi_5_awaddr,s_axi_4_awaddr,s_axi_3_awaddr,s_axi_2_awaddr,s_axi_1_awaddr,s_axi_0_awaddr};
            assign s_axi_awlen = {s_axi_9_awlen,s_axi_8_awlen,s_axi_7_awlen,s_axi_6_awlen,s_axi_5_awlen,s_axi_4_awlen,s_axi_3_awlen,s_axi_2_awlen,s_axi_1_awlen,s_axi_0_awlen};
            assign s_axi_awsize = {s_axi_9_awsize,s_axi_8_awsize,s_axi_7_awsize,s_axi_6_awsize,s_axi_5_awsize,s_axi_4_awsize,s_axi_3_awsize,s_axi_2_awsize,s_axi_1_awsize,s_axi_0_awsize};
            assign s_axi_awburst = {s_axi_9_awburst,s_axi_8_awburst,s_axi_7_awburst,s_axi_6_awburst,s_axi_5_awburst,s_axi_4_awburst,s_axi_3_awburst,s_axi_2_awburst,s_axi_1_awburst,s_axi_0_awburst};
            assign s_axi_awlock = {s_axi_9_awlock,s_axi_8_awlock,s_axi_7_awlock,s_axi_6_awlock,s_axi_5_awlock,s_axi_4_awlock,s_axi_3_awlock,s_axi_2_awlock,s_axi_1_awlock,s_axi_0_awlock};
            assign s_axi_awcache = {s_axi_9_awcache,s_axi_8_awcache,s_axi_7_awcache,s_axi_6_awcache,s_axi_5_awcache,s_axi_4_awcache,s_axi_3_awcache,s_axi_2_awcache,s_axi_1_awcache,s_axi_0_awcache};
            assign s_axi_awprot = {s_axi_9_awprot,s_axi_8_awprot,s_axi_7_awprot,s_axi_6_awprot,s_axi_5_awprot,s_axi_4_awprot,s_axi_3_awprot,s_axi_2_awprot,s_axi_1_awprot,s_axi_0_awprot};
            assign s_axi_awqos = {s_axi_9_awqos,s_axi_8_awqos,s_axi_7_awqos,s_axi_6_awqos,s_axi_5_awqos,s_axi_4_awqos,s_axi_3_awqos,s_axi_2_awqos,s_axi_1_awqos,s_axi_0_awqos};
            assign s_axi_awvalid = {s_axi_9_awvalid,s_axi_8_awvalid,s_axi_7_awvalid,s_axi_6_awvalid,s_axi_5_awvalid,s_axi_4_awvalid,s_axi_3_awvalid,s_axi_2_awvalid,s_axi_1_awvalid,s_axi_0_awvalid};
            assign {s_axi_9_awready,s_axi_8_awready,s_axi_7_awready,s_axi_6_awready,s_axi_5_awready,s_axi_4_awready,s_axi_3_awready,s_axi_2_awready,s_axi_1_awready,s_axi_0_awready} = s_axi_awready;
            assign s_axi_wdata = {s_axi_9_wdata,s_axi_8_wdata,s_axi_7_wdata,s_axi_6_wdata,s_axi_5_wdata,s_axi_4_wdata,s_axi_3_wdata,s_axi_2_wdata,s_axi_1_wdata,s_axi_0_wdata};
            assign s_axi_wstrb = {s_axi_9_wstrb,s_axi_8_wstrb,s_axi_7_wstrb,s_axi_6_wstrb,s_axi_5_wstrb,s_axi_4_wstrb,s_axi_3_wstrb,s_axi_2_wstrb,s_axi_1_wstrb,s_axi_0_wstrb};
            assign s_axi_wlast = {s_axi_9_wlast,s_axi_8_wlast,s_axi_7_wlast,s_axi_6_wlast,s_axi_5_wlast,s_axi_4_wlast,s_axi_3_wlast,s_axi_2_wlast,s_axi_1_wlast,s_axi_0_wlast};
            assign s_axi_wvalid = {s_axi_9_wvalid,s_axi_8_wvalid,s_axi_7_wvalid,s_axi_6_wvalid,s_axi_5_wvalid,s_axi_4_wvalid,s_axi_3_wvalid,s_axi_2_wvalid,s_axi_1_wvalid,s_axi_0_wvalid};
            assign {s_axi_9_wready,s_axi_8_wready,s_axi_7_wready,s_axi_6_wready,s_axi_5_wready,s_axi_4_wready,s_axi_3_wready,s_axi_2_wready,s_axi_1_wready,s_axi_0_wready} = s_axi_wready;
            assign {s_axi_9_bid,s_axi_8_bid,s_axi_7_bid,s_axi_6_bid,s_axi_5_bid,s_axi_4_bid,s_axi_3_bid,s_axi_2_bid,s_axi_1_bid,s_axi_0_bid} = s_axi_bid;
            assign {s_axi_9_bresp,s_axi_8_bresp,s_axi_7_bresp,s_axi_6_bresp,s_axi_5_bresp,s_axi_4_bresp,s_axi_3_bresp,s_axi_2_bresp,s_axi_1_bresp,s_axi_0_bresp} = s_axi_bresp;
            assign {s_axi_9_bvalid,s_axi_8_bvalid,s_axi_7_bvalid,s_axi_6_bvalid,s_axi_5_bvalid,s_axi_4_bvalid,s_axi_3_bvalid,s_axi_2_bvalid,s_axi_1_bvalid,s_axi_0_bvalid} = s_axi_bvalid;
            assign s_axi_bready = {s_axi_9_bready,s_axi_8_bready,s_axi_7_bready,s_axi_6_bready,s_axi_5_bready,s_axi_4_bready,s_axi_3_bready,s_axi_2_bready,s_axi_1_bready,s_axi_0_bready};
            assign s_axi_arid = {s_axi_9_arid,s_axi_8_arid,s_axi_7_arid,s_axi_6_arid,s_axi_5_arid,s_axi_4_arid,s_axi_3_arid,s_axi_2_arid,s_axi_1_arid,s_axi_0_arid};
            assign s_axi_araddr = {s_axi_9_araddr,s_axi_8_araddr,s_axi_7_araddr,s_axi_6_araddr,s_axi_5_araddr,s_axi_4_araddr,s_axi_3_araddr,s_axi_2_araddr,s_axi_1_araddr,s_axi_0_araddr};
            assign s_axi_arlen = {s_axi_9_arlen,s_axi_8_arlen,s_axi_7_arlen,s_axi_6_arlen,s_axi_5_arlen,s_axi_4_arlen,s_axi_3_arlen,s_axi_2_arlen,s_axi_1_arlen,s_axi_0_arlen};
            assign s_axi_arsize = {s_axi_9_arsize,s_axi_8_arsize,s_axi_7_arsize,s_axi_6_arsize,s_axi_5_arsize,s_axi_4_arsize,s_axi_3_arsize,s_axi_2_arsize,s_axi_1_arsize,s_axi_0_arsize};
            assign s_axi_arburst = {s_axi_9_arburst,s_axi_8_arburst,s_axi_7_arburst,s_axi_6_arburst,s_axi_5_arburst,s_axi_4_arburst,s_axi_3_arburst,s_axi_2_arburst,s_axi_1_arburst,s_axi_0_arburst};
            assign s_axi_arlock = {s_axi_9_arlock,s_axi_8_arlock,s_axi_7_arlock,s_axi_6_arlock,s_axi_5_arlock,s_axi_4_arlock,s_axi_3_arlock,s_axi_2_arlock,s_axi_1_arlock,s_axi_0_arlock};
            assign s_axi_arcache = {s_axi_9_arcache,s_axi_8_arcache,s_axi_7_arcache,s_axi_6_arcache,s_axi_5_arcache,s_axi_4_arcache,s_axi_3_arcache,s_axi_2_arcache,s_axi_1_arcache,s_axi_0_arcache};
            assign s_axi_arprot = {s_axi_9_arprot,s_axi_8_arprot,s_axi_7_arprot,s_axi_6_arprot,s_axi_5_arprot,s_axi_4_arprot,s_axi_3_arprot,s_axi_2_arprot,s_axi_1_arprot,s_axi_0_arprot};
            assign s_axi_arqos = {s_axi_9_arqos,s_axi_8_arqos,s_axi_7_arqos,s_axi_6_arqos,s_axi_5_arqos,s_axi_4_arqos,s_axi_3_arqos,s_axi_2_arqos,s_axi_1_arqos,s_axi_0_arqos};
            assign s_axi_arvalid = {s_axi_9_arvalid,s_axi_8_arvalid,s_axi_7_arvalid,s_axi_6_arvalid,s_axi_5_arvalid,s_axi_4_arvalid,s_axi_3_arvalid,s_axi_2_arvalid,s_axi_1_arvalid,s_axi_0_arvalid};
            assign {s_axi_9_arready,s_axi_8_arready,s_axi_7_arready,s_axi_6_arready,s_axi_5_arready,s_axi_4_arready,s_axi_3_arready,s_axi_2_arready,s_axi_1_arready,s_axi_0_arready} = s_axi_arready;
            assign {s_axi_9_rid,s_axi_8_rid,s_axi_7_rid,s_axi_6_rid,s_axi_5_rid,s_axi_4_rid,s_axi_3_rid,s_axi_2_rid,s_axi_1_rid,s_axi_0_rid} = s_axi_rid;
            assign {s_axi_9_rdata,s_axi_8_rdata,s_axi_7_rdata,s_axi_6_rdata,s_axi_5_rdata,s_axi_4_rdata,s_axi_3_rdata,s_axi_2_rdata,s_axi_1_rdata,s_axi_0_rdata} = s_axi_rdata;
            assign {s_axi_9_rresp,s_axi_8_rresp,s_axi_7_rresp,s_axi_6_rresp,s_axi_5_rresp,s_axi_4_rresp,s_axi_3_rresp,s_axi_2_rresp,s_axi_1_rresp,s_axi_0_rresp} = s_axi_rresp;
            assign {s_axi_9_rlast,s_axi_8_rlast,s_axi_7_rlast,s_axi_6_rlast,s_axi_5_rlast,s_axi_4_rlast,s_axi_3_rlast,s_axi_2_rlast,s_axi_1_rlast,s_axi_0_rlast} = s_axi_rlast;
            assign {s_axi_9_rvalid,s_axi_8_rvalid,s_axi_7_rvalid,s_axi_6_rvalid,s_axi_5_rvalid,s_axi_4_rvalid,s_axi_3_rvalid,s_axi_2_rvalid,s_axi_1_rvalid,s_axi_0_rvalid} = s_axi_rvalid;
            assign s_axi_rready = {s_axi_9_rready,s_axi_8_rready,s_axi_7_rready,s_axi_6_rready,s_axi_5_rready,s_axi_4_rready,s_axi_3_rready,s_axi_2_rready,s_axi_1_rready,s_axi_0_rready};
        end
        11: begin
            assign s_axi_awid = {s_axi_10_awid,s_axi_9_awid,s_axi_8_awid,s_axi_7_awid,s_axi_6_awid,s_axi_5_awid,s_axi_4_awid,s_axi_3_awid,s_axi_2_awid,s_axi_1_awid,s_axi_0_awid};
            assign s_axi_awaddr = {s_axi_10_awaddr,s_axi_9_awaddr,s_axi_8_awaddr,s_axi_7_awaddr,s_axi_6_awaddr,s_axi_5_awaddr,s_axi_4_awaddr,s_axi_3_awaddr,s_axi_2_awaddr,s_axi_1_awaddr,s_axi_0_awaddr};
            assign s_axi_awlen = {s_axi_10_awlen,s_axi_9_awlen,s_axi_8_awlen,s_axi_7_awlen,s_axi_6_awlen,s_axi_5_awlen,s_axi_4_awlen,s_axi_3_awlen,s_axi_2_awlen,s_axi_1_awlen,s_axi_0_awlen};
            assign s_axi_awsize = {s_axi_10_awsize,s_axi_9_awsize,s_axi_8_awsize,s_axi_7_awsize,s_axi_6_awsize,s_axi_5_awsize,s_axi_4_awsize,s_axi_3_awsize,s_axi_2_awsize,s_axi_1_awsize,s_axi_0_awsize};
            assign s_axi_awburst = {s_axi_10_awburst,s_axi_9_awburst,s_axi_8_awburst,s_axi_7_awburst,s_axi_6_awburst,s_axi_5_awburst,s_axi_4_awburst,s_axi_3_awburst,s_axi_2_awburst,s_axi_1_awburst,s_axi_0_awburst};
            assign s_axi_awlock = {s_axi_10_awlock,s_axi_9_awlock,s_axi_8_awlock,s_axi_7_awlock,s_axi_6_awlock,s_axi_5_awlock,s_axi_4_awlock,s_axi_3_awlock,s_axi_2_awlock,s_axi_1_awlock,s_axi_0_awlock};
            assign s_axi_awcache = {s_axi_10_awcache,s_axi_9_awcache,s_axi_8_awcache,s_axi_7_awcache,s_axi_6_awcache,s_axi_5_awcache,s_axi_4_awcache,s_axi_3_awcache,s_axi_2_awcache,s_axi_1_awcache,s_axi_0_awcache};
            assign s_axi_awprot = {s_axi_10_awprot,s_axi_9_awprot,s_axi_8_awprot,s_axi_7_awprot,s_axi_6_awprot,s_axi_5_awprot,s_axi_4_awprot,s_axi_3_awprot,s_axi_2_awprot,s_axi_1_awprot,s_axi_0_awprot};
            assign s_axi_awqos = {s_axi_10_awqos,s_axi_9_awqos,s_axi_8_awqos,s_axi_7_awqos,s_axi_6_awqos,s_axi_5_awqos,s_axi_4_awqos,s_axi_3_awqos,s_axi_2_awqos,s_axi_1_awqos,s_axi_0_awqos};
            assign s_axi_awvalid = {s_axi_10_awvalid,s_axi_9_awvalid,s_axi_8_awvalid,s_axi_7_awvalid,s_axi_6_awvalid,s_axi_5_awvalid,s_axi_4_awvalid,s_axi_3_awvalid,s_axi_2_awvalid,s_axi_1_awvalid,s_axi_0_awvalid};
            assign {s_axi_10_awready,s_axi_9_awready,s_axi_8_awready,s_axi_7_awready,s_axi_6_awready,s_axi_5_awready,s_axi_4_awready,s_axi_3_awready,s_axi_2_awready,s_axi_1_awready,s_axi_0_awready} = s_axi_awready;
            assign s_axi_wdata = {s_axi_10_wdata,s_axi_9_wdata,s_axi_8_wdata,s_axi_7_wdata,s_axi_6_wdata,s_axi_5_wdata,s_axi_4_wdata,s_axi_3_wdata,s_axi_2_wdata,s_axi_1_wdata,s_axi_0_wdata};
            assign s_axi_wstrb = {s_axi_10_wstrb,s_axi_9_wstrb,s_axi_8_wstrb,s_axi_7_wstrb,s_axi_6_wstrb,s_axi_5_wstrb,s_axi_4_wstrb,s_axi_3_wstrb,s_axi_2_wstrb,s_axi_1_wstrb,s_axi_0_wstrb};
            assign s_axi_wlast = {s_axi_10_wlast,s_axi_9_wlast,s_axi_8_wlast,s_axi_7_wlast,s_axi_6_wlast,s_axi_5_wlast,s_axi_4_wlast,s_axi_3_wlast,s_axi_2_wlast,s_axi_1_wlast,s_axi_0_wlast};
            assign s_axi_wvalid = {s_axi_10_wvalid,s_axi_9_wvalid,s_axi_8_wvalid,s_axi_7_wvalid,s_axi_6_wvalid,s_axi_5_wvalid,s_axi_4_wvalid,s_axi_3_wvalid,s_axi_2_wvalid,s_axi_1_wvalid,s_axi_0_wvalid};
            assign {s_axi_10_wready,s_axi_9_wready,s_axi_8_wready,s_axi_7_wready,s_axi_6_wready,s_axi_5_wready,s_axi_4_wready,s_axi_3_wready,s_axi_2_wready,s_axi_1_wready,s_axi_0_wready} = s_axi_wready;
            assign {s_axi_10_bid,s_axi_9_bid,s_axi_8_bid,s_axi_7_bid,s_axi_6_bid,s_axi_5_bid,s_axi_4_bid,s_axi_3_bid,s_axi_2_bid,s_axi_1_bid,s_axi_0_bid} = s_axi_bid;
            assign {s_axi_10_bresp,s_axi_9_bresp,s_axi_8_bresp,s_axi_7_bresp,s_axi_6_bresp,s_axi_5_bresp,s_axi_4_bresp,s_axi_3_bresp,s_axi_2_bresp,s_axi_1_bresp,s_axi_0_bresp} = s_axi_bresp;
            assign {s_axi_10_bvalid,s_axi_9_bvalid,s_axi_8_bvalid,s_axi_7_bvalid,s_axi_6_bvalid,s_axi_5_bvalid,s_axi_4_bvalid,s_axi_3_bvalid,s_axi_2_bvalid,s_axi_1_bvalid,s_axi_0_bvalid} = s_axi_bvalid;
            assign s_axi_bready = {s_axi_10_bready,s_axi_9_bready,s_axi_8_bready,s_axi_7_bready,s_axi_6_bready,s_axi_5_bready,s_axi_4_bready,s_axi_3_bready,s_axi_2_bready,s_axi_1_bready,s_axi_0_bready};
            assign s_axi_arid = {s_axi_10_arid,s_axi_9_arid,s_axi_8_arid,s_axi_7_arid,s_axi_6_arid,s_axi_5_arid,s_axi_4_arid,s_axi_3_arid,s_axi_2_arid,s_axi_1_arid,s_axi_0_arid};
            assign s_axi_araddr = {s_axi_10_araddr,s_axi_9_araddr,s_axi_8_araddr,s_axi_7_araddr,s_axi_6_araddr,s_axi_5_araddr,s_axi_4_araddr,s_axi_3_araddr,s_axi_2_araddr,s_axi_1_araddr,s_axi_0_araddr};
            assign s_axi_arlen = {s_axi_10_arlen,s_axi_9_arlen,s_axi_8_arlen,s_axi_7_arlen,s_axi_6_arlen,s_axi_5_arlen,s_axi_4_arlen,s_axi_3_arlen,s_axi_2_arlen,s_axi_1_arlen,s_axi_0_arlen};
            assign s_axi_arsize = {s_axi_10_arsize,s_axi_9_arsize,s_axi_8_arsize,s_axi_7_arsize,s_axi_6_arsize,s_axi_5_arsize,s_axi_4_arsize,s_axi_3_arsize,s_axi_2_arsize,s_axi_1_arsize,s_axi_0_arsize};
            assign s_axi_arburst = {s_axi_10_arburst,s_axi_9_arburst,s_axi_8_arburst,s_axi_7_arburst,s_axi_6_arburst,s_axi_5_arburst,s_axi_4_arburst,s_axi_3_arburst,s_axi_2_arburst,s_axi_1_arburst,s_axi_0_arburst};
            assign s_axi_arlock = {s_axi_10_arlock,s_axi_9_arlock,s_axi_8_arlock,s_axi_7_arlock,s_axi_6_arlock,s_axi_5_arlock,s_axi_4_arlock,s_axi_3_arlock,s_axi_2_arlock,s_axi_1_arlock,s_axi_0_arlock};
            assign s_axi_arcache = {s_axi_10_arcache,s_axi_9_arcache,s_axi_8_arcache,s_axi_7_arcache,s_axi_6_arcache,s_axi_5_arcache,s_axi_4_arcache,s_axi_3_arcache,s_axi_2_arcache,s_axi_1_arcache,s_axi_0_arcache};
            assign s_axi_arprot = {s_axi_10_arprot,s_axi_9_arprot,s_axi_8_arprot,s_axi_7_arprot,s_axi_6_arprot,s_axi_5_arprot,s_axi_4_arprot,s_axi_3_arprot,s_axi_2_arprot,s_axi_1_arprot,s_axi_0_arprot};
            assign s_axi_arqos = {s_axi_10_arqos,s_axi_9_arqos,s_axi_8_arqos,s_axi_7_arqos,s_axi_6_arqos,s_axi_5_arqos,s_axi_4_arqos,s_axi_3_arqos,s_axi_2_arqos,s_axi_1_arqos,s_axi_0_arqos};
            assign s_axi_arvalid = {s_axi_10_arvalid,s_axi_9_arvalid,s_axi_8_arvalid,s_axi_7_arvalid,s_axi_6_arvalid,s_axi_5_arvalid,s_axi_4_arvalid,s_axi_3_arvalid,s_axi_2_arvalid,s_axi_1_arvalid,s_axi_0_arvalid};
            assign {s_axi_10_arready,s_axi_9_arready,s_axi_8_arready,s_axi_7_arready,s_axi_6_arready,s_axi_5_arready,s_axi_4_arready,s_axi_3_arready,s_axi_2_arready,s_axi_1_arready,s_axi_0_arready} = s_axi_arready;
            assign {s_axi_10_rid,s_axi_9_rid,s_axi_8_rid,s_axi_7_rid,s_axi_6_rid,s_axi_5_rid,s_axi_4_rid,s_axi_3_rid,s_axi_2_rid,s_axi_1_rid,s_axi_0_rid} = s_axi_rid;
            assign {s_axi_10_rdata,s_axi_9_rdata,s_axi_8_rdata,s_axi_7_rdata,s_axi_6_rdata,s_axi_5_rdata,s_axi_4_rdata,s_axi_3_rdata,s_axi_2_rdata,s_axi_1_rdata,s_axi_0_rdata} = s_axi_rdata;
            assign {s_axi_10_rresp,s_axi_9_rresp,s_axi_8_rresp,s_axi_7_rresp,s_axi_6_rresp,s_axi_5_rresp,s_axi_4_rresp,s_axi_3_rresp,s_axi_2_rresp,s_axi_1_rresp,s_axi_0_rresp} = s_axi_rresp;
            assign {s_axi_10_rlast,s_axi_9_rlast,s_axi_8_rlast,s_axi_7_rlast,s_axi_6_rlast,s_axi_5_rlast,s_axi_4_rlast,s_axi_3_rlast,s_axi_2_rlast,s_axi_1_rlast,s_axi_0_rlast} = s_axi_rlast;
            assign {s_axi_10_rvalid,s_axi_9_rvalid,s_axi_8_rvalid,s_axi_7_rvalid,s_axi_6_rvalid,s_axi_5_rvalid,s_axi_4_rvalid,s_axi_3_rvalid,s_axi_2_rvalid,s_axi_1_rvalid,s_axi_0_rvalid} = s_axi_rvalid;
            assign s_axi_rready = {s_axi_10_rready,s_axi_9_rready,s_axi_8_rready,s_axi_7_rready,s_axi_6_rready,s_axi_5_rready,s_axi_4_rready,s_axi_3_rready,s_axi_2_rready,s_axi_1_rready,s_axi_0_rready};
        end
        12: begin
            assign s_axi_awid = {s_axi_11_awid,s_axi_10_awid,s_axi_9_awid,s_axi_8_awid,s_axi_7_awid,s_axi_6_awid,s_axi_5_awid,s_axi_4_awid,s_axi_3_awid,s_axi_2_awid,s_axi_1_awid,s_axi_0_awid};
            assign s_axi_awaddr = {s_axi_11_awaddr,s_axi_10_awaddr,s_axi_9_awaddr,s_axi_8_awaddr,s_axi_7_awaddr,s_axi_6_awaddr,s_axi_5_awaddr,s_axi_4_awaddr,s_axi_3_awaddr,s_axi_2_awaddr,s_axi_1_awaddr,s_axi_0_awaddr};
            assign s_axi_awlen = {s_axi_11_awlen,s_axi_10_awlen,s_axi_9_awlen,s_axi_8_awlen,s_axi_7_awlen,s_axi_6_awlen,s_axi_5_awlen,s_axi_4_awlen,s_axi_3_awlen,s_axi_2_awlen,s_axi_1_awlen,s_axi_0_awlen};
            assign s_axi_awsize = {s_axi_11_awsize,s_axi_10_awsize,s_axi_9_awsize,s_axi_8_awsize,s_axi_7_awsize,s_axi_6_awsize,s_axi_5_awsize,s_axi_4_awsize,s_axi_3_awsize,s_axi_2_awsize,s_axi_1_awsize,s_axi_0_awsize};
            assign s_axi_awburst = {s_axi_11_awburst,s_axi_10_awburst,s_axi_9_awburst,s_axi_8_awburst,s_axi_7_awburst,s_axi_6_awburst,s_axi_5_awburst,s_axi_4_awburst,s_axi_3_awburst,s_axi_2_awburst,s_axi_1_awburst,s_axi_0_awburst};
            assign s_axi_awlock = {s_axi_11_awlock,s_axi_10_awlock,s_axi_9_awlock,s_axi_8_awlock,s_axi_7_awlock,s_axi_6_awlock,s_axi_5_awlock,s_axi_4_awlock,s_axi_3_awlock,s_axi_2_awlock,s_axi_1_awlock,s_axi_0_awlock};
            assign s_axi_awcache = {s_axi_11_awcache,s_axi_10_awcache,s_axi_9_awcache,s_axi_8_awcache,s_axi_7_awcache,s_axi_6_awcache,s_axi_5_awcache,s_axi_4_awcache,s_axi_3_awcache,s_axi_2_awcache,s_axi_1_awcache,s_axi_0_awcache};
            assign s_axi_awprot = {s_axi_11_awprot,s_axi_10_awprot,s_axi_9_awprot,s_axi_8_awprot,s_axi_7_awprot,s_axi_6_awprot,s_axi_5_awprot,s_axi_4_awprot,s_axi_3_awprot,s_axi_2_awprot,s_axi_1_awprot,s_axi_0_awprot};
            assign s_axi_awqos = {s_axi_11_awqos,s_axi_10_awqos,s_axi_9_awqos,s_axi_8_awqos,s_axi_7_awqos,s_axi_6_awqos,s_axi_5_awqos,s_axi_4_awqos,s_axi_3_awqos,s_axi_2_awqos,s_axi_1_awqos,s_axi_0_awqos};
            assign s_axi_awvalid = {s_axi_11_awvalid,s_axi_10_awvalid,s_axi_9_awvalid,s_axi_8_awvalid,s_axi_7_awvalid,s_axi_6_awvalid,s_axi_5_awvalid,s_axi_4_awvalid,s_axi_3_awvalid,s_axi_2_awvalid,s_axi_1_awvalid,s_axi_0_awvalid};
            assign {s_axi_11_awready,s_axi_10_awready,s_axi_9_awready,s_axi_8_awready,s_axi_7_awready,s_axi_6_awready,s_axi_5_awready,s_axi_4_awready,s_axi_3_awready,s_axi_2_awready,s_axi_1_awready,s_axi_0_awready} = s_axi_awready;
            assign s_axi_wdata = {s_axi_11_wdata,s_axi_10_wdata,s_axi_9_wdata,s_axi_8_wdata,s_axi_7_wdata,s_axi_6_wdata,s_axi_5_wdata,s_axi_4_wdata,s_axi_3_wdata,s_axi_2_wdata,s_axi_1_wdata,s_axi_0_wdata};
            assign s_axi_wstrb = {s_axi_11_wstrb,s_axi_10_wstrb,s_axi_9_wstrb,s_axi_8_wstrb,s_axi_7_wstrb,s_axi_6_wstrb,s_axi_5_wstrb,s_axi_4_wstrb,s_axi_3_wstrb,s_axi_2_wstrb,s_axi_1_wstrb,s_axi_0_wstrb};
            assign s_axi_wlast = {s_axi_11_wlast,s_axi_10_wlast,s_axi_9_wlast,s_axi_8_wlast,s_axi_7_wlast,s_axi_6_wlast,s_axi_5_wlast,s_axi_4_wlast,s_axi_3_wlast,s_axi_2_wlast,s_axi_1_wlast,s_axi_0_wlast};
            assign s_axi_wvalid = {s_axi_11_wvalid,s_axi_10_wvalid,s_axi_9_wvalid,s_axi_8_wvalid,s_axi_7_wvalid,s_axi_6_wvalid,s_axi_5_wvalid,s_axi_4_wvalid,s_axi_3_wvalid,s_axi_2_wvalid,s_axi_1_wvalid,s_axi_0_wvalid};
            assign {s_axi_11_wready,s_axi_10_wready,s_axi_9_wready,s_axi_8_wready,s_axi_7_wready,s_axi_6_wready,s_axi_5_wready,s_axi_4_wready,s_axi_3_wready,s_axi_2_wready,s_axi_1_wready,s_axi_0_wready} = s_axi_wready;
            assign {s_axi_11_bid,s_axi_10_bid,s_axi_9_bid,s_axi_8_bid,s_axi_7_bid,s_axi_6_bid,s_axi_5_bid,s_axi_4_bid,s_axi_3_bid,s_axi_2_bid,s_axi_1_bid,s_axi_0_bid} = s_axi_bid;
            assign {s_axi_11_bresp,s_axi_10_bresp,s_axi_9_bresp,s_axi_8_bresp,s_axi_7_bresp,s_axi_6_bresp,s_axi_5_bresp,s_axi_4_bresp,s_axi_3_bresp,s_axi_2_bresp,s_axi_1_bresp,s_axi_0_bresp} = s_axi_bresp;
            assign {s_axi_11_bvalid,s_axi_10_bvalid,s_axi_9_bvalid,s_axi_8_bvalid,s_axi_7_bvalid,s_axi_6_bvalid,s_axi_5_bvalid,s_axi_4_bvalid,s_axi_3_bvalid,s_axi_2_bvalid,s_axi_1_bvalid,s_axi_0_bvalid} = s_axi_bvalid;
            assign s_axi_bready = {s_axi_11_bready,s_axi_10_bready,s_axi_9_bready,s_axi_8_bready,s_axi_7_bready,s_axi_6_bready,s_axi_5_bready,s_axi_4_bready,s_axi_3_bready,s_axi_2_bready,s_axi_1_bready,s_axi_0_bready};
            assign s_axi_arid = {s_axi_11_arid,s_axi_10_arid,s_axi_9_arid,s_axi_8_arid,s_axi_7_arid,s_axi_6_arid,s_axi_5_arid,s_axi_4_arid,s_axi_3_arid,s_axi_2_arid,s_axi_1_arid,s_axi_0_arid};
            assign s_axi_araddr = {s_axi_11_araddr,s_axi_10_araddr,s_axi_9_araddr,s_axi_8_araddr,s_axi_7_araddr,s_axi_6_araddr,s_axi_5_araddr,s_axi_4_araddr,s_axi_3_araddr,s_axi_2_araddr,s_axi_1_araddr,s_axi_0_araddr};
            assign s_axi_arlen = {s_axi_11_arlen,s_axi_10_arlen,s_axi_9_arlen,s_axi_8_arlen,s_axi_7_arlen,s_axi_6_arlen,s_axi_5_arlen,s_axi_4_arlen,s_axi_3_arlen,s_axi_2_arlen,s_axi_1_arlen,s_axi_0_arlen};
            assign s_axi_arsize = {s_axi_11_arsize,s_axi_10_arsize,s_axi_9_arsize,s_axi_8_arsize,s_axi_7_arsize,s_axi_6_arsize,s_axi_5_arsize,s_axi_4_arsize,s_axi_3_arsize,s_axi_2_arsize,s_axi_1_arsize,s_axi_0_arsize};
            assign s_axi_arburst = {s_axi_11_arburst,s_axi_10_arburst,s_axi_9_arburst,s_axi_8_arburst,s_axi_7_arburst,s_axi_6_arburst,s_axi_5_arburst,s_axi_4_arburst,s_axi_3_arburst,s_axi_2_arburst,s_axi_1_arburst,s_axi_0_arburst};
            assign s_axi_arlock = {s_axi_11_arlock,s_axi_10_arlock,s_axi_9_arlock,s_axi_8_arlock,s_axi_7_arlock,s_axi_6_arlock,s_axi_5_arlock,s_axi_4_arlock,s_axi_3_arlock,s_axi_2_arlock,s_axi_1_arlock,s_axi_0_arlock};
            assign s_axi_arcache = {s_axi_11_arcache,s_axi_10_arcache,s_axi_9_arcache,s_axi_8_arcache,s_axi_7_arcache,s_axi_6_arcache,s_axi_5_arcache,s_axi_4_arcache,s_axi_3_arcache,s_axi_2_arcache,s_axi_1_arcache,s_axi_0_arcache};
            assign s_axi_arprot = {s_axi_11_arprot,s_axi_10_arprot,s_axi_9_arprot,s_axi_8_arprot,s_axi_7_arprot,s_axi_6_arprot,s_axi_5_arprot,s_axi_4_arprot,s_axi_3_arprot,s_axi_2_arprot,s_axi_1_arprot,s_axi_0_arprot};
            assign s_axi_arqos = {s_axi_11_arqos,s_axi_10_arqos,s_axi_9_arqos,s_axi_8_arqos,s_axi_7_arqos,s_axi_6_arqos,s_axi_5_arqos,s_axi_4_arqos,s_axi_3_arqos,s_axi_2_arqos,s_axi_1_arqos,s_axi_0_arqos};
            assign s_axi_arvalid = {s_axi_11_arvalid,s_axi_10_arvalid,s_axi_9_arvalid,s_axi_8_arvalid,s_axi_7_arvalid,s_axi_6_arvalid,s_axi_5_arvalid,s_axi_4_arvalid,s_axi_3_arvalid,s_axi_2_arvalid,s_axi_1_arvalid,s_axi_0_arvalid};
            assign {s_axi_11_arready,s_axi_10_arready,s_axi_9_arready,s_axi_8_arready,s_axi_7_arready,s_axi_6_arready,s_axi_5_arready,s_axi_4_arready,s_axi_3_arready,s_axi_2_arready,s_axi_1_arready,s_axi_0_arready} = s_axi_arready;
            assign {s_axi_11_rid,s_axi_10_rid,s_axi_9_rid,s_axi_8_rid,s_axi_7_rid,s_axi_6_rid,s_axi_5_rid,s_axi_4_rid,s_axi_3_rid,s_axi_2_rid,s_axi_1_rid,s_axi_0_rid} = s_axi_rid;
            assign {s_axi_11_rdata,s_axi_10_rdata,s_axi_9_rdata,s_axi_8_rdata,s_axi_7_rdata,s_axi_6_rdata,s_axi_5_rdata,s_axi_4_rdata,s_axi_3_rdata,s_axi_2_rdata,s_axi_1_rdata,s_axi_0_rdata} = s_axi_rdata;
            assign {s_axi_11_rresp,s_axi_10_rresp,s_axi_9_rresp,s_axi_8_rresp,s_axi_7_rresp,s_axi_6_rresp,s_axi_5_rresp,s_axi_4_rresp,s_axi_3_rresp,s_axi_2_rresp,s_axi_1_rresp,s_axi_0_rresp} = s_axi_rresp;
            assign {s_axi_11_rlast,s_axi_10_rlast,s_axi_9_rlast,s_axi_8_rlast,s_axi_7_rlast,s_axi_6_rlast,s_axi_5_rlast,s_axi_4_rlast,s_axi_3_rlast,s_axi_2_rlast,s_axi_1_rlast,s_axi_0_rlast} = s_axi_rlast;
            assign {s_axi_11_rvalid,s_axi_10_rvalid,s_axi_9_rvalid,s_axi_8_rvalid,s_axi_7_rvalid,s_axi_6_rvalid,s_axi_5_rvalid,s_axi_4_rvalid,s_axi_3_rvalid,s_axi_2_rvalid,s_axi_1_rvalid,s_axi_0_rvalid} = s_axi_rvalid;
            assign s_axi_rready = {s_axi_11_rready,s_axi_10_rready,s_axi_9_rready,s_axi_8_rready,s_axi_7_rready,s_axi_6_rready,s_axi_5_rready,s_axi_4_rready,s_axi_3_rready,s_axi_2_rready,s_axi_1_rready,s_axi_0_rready};
        end
        13: begin
            assign s_axi_awid = {s_axi_12_awid,s_axi_11_awid,s_axi_10_awid,s_axi_9_awid,s_axi_8_awid,s_axi_7_awid,s_axi_6_awid,s_axi_5_awid,s_axi_4_awid,s_axi_3_awid,s_axi_2_awid,s_axi_1_awid,s_axi_0_awid};
            assign s_axi_awaddr = {s_axi_12_awaddr,s_axi_11_awaddr,s_axi_10_awaddr,s_axi_9_awaddr,s_axi_8_awaddr,s_axi_7_awaddr,s_axi_6_awaddr,s_axi_5_awaddr,s_axi_4_awaddr,s_axi_3_awaddr,s_axi_2_awaddr,s_axi_1_awaddr,s_axi_0_awaddr};
            assign s_axi_awlen = {s_axi_12_awlen,s_axi_11_awlen,s_axi_10_awlen,s_axi_9_awlen,s_axi_8_awlen,s_axi_7_awlen,s_axi_6_awlen,s_axi_5_awlen,s_axi_4_awlen,s_axi_3_awlen,s_axi_2_awlen,s_axi_1_awlen,s_axi_0_awlen};
            assign s_axi_awsize = {s_axi_12_awsize,s_axi_11_awsize,s_axi_10_awsize,s_axi_9_awsize,s_axi_8_awsize,s_axi_7_awsize,s_axi_6_awsize,s_axi_5_awsize,s_axi_4_awsize,s_axi_3_awsize,s_axi_2_awsize,s_axi_1_awsize,s_axi_0_awsize};
            assign s_axi_awburst = {s_axi_12_awburst,s_axi_11_awburst,s_axi_10_awburst,s_axi_9_awburst,s_axi_8_awburst,s_axi_7_awburst,s_axi_6_awburst,s_axi_5_awburst,s_axi_4_awburst,s_axi_3_awburst,s_axi_2_awburst,s_axi_1_awburst,s_axi_0_awburst};
            assign s_axi_awlock = {s_axi_12_awlock,s_axi_11_awlock,s_axi_10_awlock,s_axi_9_awlock,s_axi_8_awlock,s_axi_7_awlock,s_axi_6_awlock,s_axi_5_awlock,s_axi_4_awlock,s_axi_3_awlock,s_axi_2_awlock,s_axi_1_awlock,s_axi_0_awlock};
            assign s_axi_awcache = {s_axi_12_awcache,s_axi_11_awcache,s_axi_10_awcache,s_axi_9_awcache,s_axi_8_awcache,s_axi_7_awcache,s_axi_6_awcache,s_axi_5_awcache,s_axi_4_awcache,s_axi_3_awcache,s_axi_2_awcache,s_axi_1_awcache,s_axi_0_awcache};
            assign s_axi_awprot = {s_axi_12_awprot,s_axi_11_awprot,s_axi_10_awprot,s_axi_9_awprot,s_axi_8_awprot,s_axi_7_awprot,s_axi_6_awprot,s_axi_5_awprot,s_axi_4_awprot,s_axi_3_awprot,s_axi_2_awprot,s_axi_1_awprot,s_axi_0_awprot};
            assign s_axi_awqos = {s_axi_12_awqos,s_axi_11_awqos,s_axi_10_awqos,s_axi_9_awqos,s_axi_8_awqos,s_axi_7_awqos,s_axi_6_awqos,s_axi_5_awqos,s_axi_4_awqos,s_axi_3_awqos,s_axi_2_awqos,s_axi_1_awqos,s_axi_0_awqos};
            assign s_axi_awvalid = {s_axi_12_awvalid,s_axi_11_awvalid,s_axi_10_awvalid,s_axi_9_awvalid,s_axi_8_awvalid,s_axi_7_awvalid,s_axi_6_awvalid,s_axi_5_awvalid,s_axi_4_awvalid,s_axi_3_awvalid,s_axi_2_awvalid,s_axi_1_awvalid,s_axi_0_awvalid};
            assign {s_axi_12_awready,s_axi_11_awready,s_axi_10_awready,s_axi_9_awready,s_axi_8_awready,s_axi_7_awready,s_axi_6_awready,s_axi_5_awready,s_axi_4_awready,s_axi_3_awready,s_axi_2_awready,s_axi_1_awready,s_axi_0_awready} = s_axi_awready;
            assign s_axi_wdata = {s_axi_12_wdata,s_axi_11_wdata,s_axi_10_wdata,s_axi_9_wdata,s_axi_8_wdata,s_axi_7_wdata,s_axi_6_wdata,s_axi_5_wdata,s_axi_4_wdata,s_axi_3_wdata,s_axi_2_wdata,s_axi_1_wdata,s_axi_0_wdata};
            assign s_axi_wstrb = {s_axi_12_wstrb,s_axi_11_wstrb,s_axi_10_wstrb,s_axi_9_wstrb,s_axi_8_wstrb,s_axi_7_wstrb,s_axi_6_wstrb,s_axi_5_wstrb,s_axi_4_wstrb,s_axi_3_wstrb,s_axi_2_wstrb,s_axi_1_wstrb,s_axi_0_wstrb};
            assign s_axi_wlast = {s_axi_12_wlast,s_axi_11_wlast,s_axi_10_wlast,s_axi_9_wlast,s_axi_8_wlast,s_axi_7_wlast,s_axi_6_wlast,s_axi_5_wlast,s_axi_4_wlast,s_axi_3_wlast,s_axi_2_wlast,s_axi_1_wlast,s_axi_0_wlast};
            assign s_axi_wvalid = {s_axi_12_wvalid,s_axi_11_wvalid,s_axi_10_wvalid,s_axi_9_wvalid,s_axi_8_wvalid,s_axi_7_wvalid,s_axi_6_wvalid,s_axi_5_wvalid,s_axi_4_wvalid,s_axi_3_wvalid,s_axi_2_wvalid,s_axi_1_wvalid,s_axi_0_wvalid};
            assign {s_axi_12_wready,s_axi_11_wready,s_axi_10_wready,s_axi_9_wready,s_axi_8_wready,s_axi_7_wready,s_axi_6_wready,s_axi_5_wready,s_axi_4_wready,s_axi_3_wready,s_axi_2_wready,s_axi_1_wready,s_axi_0_wready} = s_axi_wready;
            assign {s_axi_12_bid,s_axi_11_bid,s_axi_10_bid,s_axi_9_bid,s_axi_8_bid,s_axi_7_bid,s_axi_6_bid,s_axi_5_bid,s_axi_4_bid,s_axi_3_bid,s_axi_2_bid,s_axi_1_bid,s_axi_0_bid} = s_axi_bid;
            assign {s_axi_12_bresp,s_axi_11_bresp,s_axi_10_bresp,s_axi_9_bresp,s_axi_8_bresp,s_axi_7_bresp,s_axi_6_bresp,s_axi_5_bresp,s_axi_4_bresp,s_axi_3_bresp,s_axi_2_bresp,s_axi_1_bresp,s_axi_0_bresp} = s_axi_bresp;
            assign {s_axi_12_bvalid,s_axi_11_bvalid,s_axi_10_bvalid,s_axi_9_bvalid,s_axi_8_bvalid,s_axi_7_bvalid,s_axi_6_bvalid,s_axi_5_bvalid,s_axi_4_bvalid,s_axi_3_bvalid,s_axi_2_bvalid,s_axi_1_bvalid,s_axi_0_bvalid} = s_axi_bvalid;
            assign s_axi_bready = {s_axi_12_bready,s_axi_11_bready,s_axi_10_bready,s_axi_9_bready,s_axi_8_bready,s_axi_7_bready,s_axi_6_bready,s_axi_5_bready,s_axi_4_bready,s_axi_3_bready,s_axi_2_bready,s_axi_1_bready,s_axi_0_bready};
            assign s_axi_arid = {s_axi_12_arid,s_axi_11_arid,s_axi_10_arid,s_axi_9_arid,s_axi_8_arid,s_axi_7_arid,s_axi_6_arid,s_axi_5_arid,s_axi_4_arid,s_axi_3_arid,s_axi_2_arid,s_axi_1_arid,s_axi_0_arid};
            assign s_axi_araddr = {s_axi_12_araddr,s_axi_11_araddr,s_axi_10_araddr,s_axi_9_araddr,s_axi_8_araddr,s_axi_7_araddr,s_axi_6_araddr,s_axi_5_araddr,s_axi_4_araddr,s_axi_3_araddr,s_axi_2_araddr,s_axi_1_araddr,s_axi_0_araddr};
            assign s_axi_arlen = {s_axi_12_arlen,s_axi_11_arlen,s_axi_10_arlen,s_axi_9_arlen,s_axi_8_arlen,s_axi_7_arlen,s_axi_6_arlen,s_axi_5_arlen,s_axi_4_arlen,s_axi_3_arlen,s_axi_2_arlen,s_axi_1_arlen,s_axi_0_arlen};
            assign s_axi_arsize = {s_axi_12_arsize,s_axi_11_arsize,s_axi_10_arsize,s_axi_9_arsize,s_axi_8_arsize,s_axi_7_arsize,s_axi_6_arsize,s_axi_5_arsize,s_axi_4_arsize,s_axi_3_arsize,s_axi_2_arsize,s_axi_1_arsize,s_axi_0_arsize};
            assign s_axi_arburst = {s_axi_12_arburst,s_axi_11_arburst,s_axi_10_arburst,s_axi_9_arburst,s_axi_8_arburst,s_axi_7_arburst,s_axi_6_arburst,s_axi_5_arburst,s_axi_4_arburst,s_axi_3_arburst,s_axi_2_arburst,s_axi_1_arburst,s_axi_0_arburst};
            assign s_axi_arlock = {s_axi_12_arlock,s_axi_11_arlock,s_axi_10_arlock,s_axi_9_arlock,s_axi_8_arlock,s_axi_7_arlock,s_axi_6_arlock,s_axi_5_arlock,s_axi_4_arlock,s_axi_3_arlock,s_axi_2_arlock,s_axi_1_arlock,s_axi_0_arlock};
            assign s_axi_arcache = {s_axi_12_arcache,s_axi_11_arcache,s_axi_10_arcache,s_axi_9_arcache,s_axi_8_arcache,s_axi_7_arcache,s_axi_6_arcache,s_axi_5_arcache,s_axi_4_arcache,s_axi_3_arcache,s_axi_2_arcache,s_axi_1_arcache,s_axi_0_arcache};
            assign s_axi_arprot = {s_axi_12_arprot,s_axi_11_arprot,s_axi_10_arprot,s_axi_9_arprot,s_axi_8_arprot,s_axi_7_arprot,s_axi_6_arprot,s_axi_5_arprot,s_axi_4_arprot,s_axi_3_arprot,s_axi_2_arprot,s_axi_1_arprot,s_axi_0_arprot};
            assign s_axi_arqos = {s_axi_12_arqos,s_axi_11_arqos,s_axi_10_arqos,s_axi_9_arqos,s_axi_8_arqos,s_axi_7_arqos,s_axi_6_arqos,s_axi_5_arqos,s_axi_4_arqos,s_axi_3_arqos,s_axi_2_arqos,s_axi_1_arqos,s_axi_0_arqos};
            assign {s_axi_12_arvalid,s_axi_11_arvalid,s_axi_10_arvalid,s_axi_9_arvalid,s_axi_8_arvalid,s_axi_7_arvalid,s_axi_6_arvalid,s_axi_5_arvalid,s_axi_4_arvalid,s_axi_3_arvalid,s_axi_2_arvalid,s_axi_1_arvalid,s_axi_0_arvalid} = s_axi_arvalid;
            assign {s_axi_12_arready,s_axi_11_arready,s_axi_10_arready,s_axi_9_arready,s_axi_8_arready,s_axi_7_arready,s_axi_6_arready,s_axi_5_arready,s_axi_4_arready,s_axi_3_arready,s_axi_2_arready,s_axi_1_arready,s_axi_0_arready} = s_axi_arready;
            assign {s_axi_12_rid,s_axi_11_rid,s_axi_10_rid,s_axi_9_rid,s_axi_8_rid,s_axi_7_rid,s_axi_6_rid,s_axi_5_rid,s_axi_4_rid,s_axi_3_rid,s_axi_2_rid,s_axi_1_rid,s_axi_0_rid} = s_axi_rid;
            assign {s_axi_12_rdata,s_axi_11_rdata,s_axi_10_rdata,s_axi_9_rdata,s_axi_8_rdata,s_axi_7_rdata,s_axi_6_rdata,s_axi_5_rdata,s_axi_4_rdata,s_axi_3_rdata,s_axi_2_rdata,s_axi_1_rdata,s_axi_0_rdata} = s_axi_rdata;
            assign {s_axi_12_rresp,s_axi_11_rresp,s_axi_10_rresp,s_axi_9_rresp,s_axi_8_rresp,s_axi_7_rresp,s_axi_6_rresp,s_axi_5_rresp,s_axi_4_rresp,s_axi_3_rresp,s_axi_2_rresp,s_axi_1_rresp,s_axi_0_rresp} = s_axi_rresp;
            assign {s_axi_12_rlast,s_axi_11_rlast,s_axi_10_rlast,s_axi_9_rlast,s_axi_8_rlast,s_axi_7_rlast,s_axi_6_rlast,s_axi_5_rlast,s_axi_4_rlast,s_axi_3_rlast,s_axi_2_rlast,s_axi_1_rlast,s_axi_0_rlast} = s_axi_rlast;
            assign {s_axi_12_rvalid,s_axi_11_rvalid,s_axi_10_rvalid,s_axi_9_rvalid,s_axi_8_rvalid,s_axi_7_rvalid,s_axi_6_rvalid,s_axi_5_rvalid,s_axi_4_rvalid,s_axi_3_rvalid,s_axi_2_rvalid,s_axi_1_rvalid,s_axi_0_rvalid} = s_axi_rvalid;
            assign s_axi_rready = {s_axi_12_rready,s_axi_11_rready,s_axi_10_rready,s_axi_9_rready,s_axi_8_rready,s_axi_7_rready,s_axi_6_rready,s_axi_5_rready,s_axi_4_rready,s_axi_3_rready,s_axi_2_rready,s_axi_1_rready,s_axi_0_rready};
        end
        14: begin
            assign s_axi_awid = {s_axi_13_awid,s_axi_12_awid,s_axi_11_awid,s_axi_10_awid,s_axi_9_awid,s_axi_8_awid,s_axi_7_awid,s_axi_6_awid,s_axi_5_awid,s_axi_4_awid,s_axi_3_awid,s_axi_2_awid,s_axi_1_awid,s_axi_0_awid};
            assign s_axi_awaddr = {s_axi_13_awaddr,s_axi_12_awaddr,s_axi_11_awaddr,s_axi_10_awaddr,s_axi_9_awaddr,s_axi_8_awaddr,s_axi_7_awaddr,s_axi_6_awaddr,s_axi_5_awaddr,s_axi_4_awaddr,s_axi_3_awaddr,s_axi_2_awaddr,s_axi_1_awaddr,s_axi_0_awaddr};
            assign s_axi_awlen = {s_axi_13_awlen,s_axi_12_awlen,s_axi_11_awlen,s_axi_10_awlen,s_axi_9_awlen,s_axi_8_awlen,s_axi_7_awlen,s_axi_6_awlen,s_axi_5_awlen,s_axi_4_awlen,s_axi_3_awlen,s_axi_2_awlen,s_axi_1_awlen,s_axi_0_awlen};
            assign s_axi_awsize = {s_axi_13_awsize,s_axi_12_awsize,s_axi_11_awsize,s_axi_10_awsize,s_axi_9_awsize,s_axi_8_awsize,s_axi_7_awsize,s_axi_6_awsize,s_axi_5_awsize,s_axi_4_awsize,s_axi_3_awsize,s_axi_2_awsize,s_axi_1_awsize,s_axi_0_awsize};
            assign s_axi_awburst = {s_axi_13_awburst,s_axi_12_awburst,s_axi_11_awburst,s_axi_10_awburst,s_axi_9_awburst,s_axi_8_awburst,s_axi_7_awburst,s_axi_6_awburst,s_axi_5_awburst,s_axi_4_awburst,s_axi_3_awburst,s_axi_2_awburst,s_axi_1_awburst,s_axi_0_awburst};
            assign s_axi_awlock = {s_axi_13_awlock,s_axi_12_awlock,s_axi_11_awlock,s_axi_10_awlock,s_axi_9_awlock,s_axi_8_awlock,s_axi_7_awlock,s_axi_6_awlock,s_axi_5_awlock,s_axi_4_awlock,s_axi_3_awlock,s_axi_2_awlock,s_axi_1_awlock,s_axi_0_awlock};
            assign s_axi_awcache = {s_axi_13_awcache,s_axi_12_awcache,s_axi_11_awcache,s_axi_10_awcache,s_axi_9_awcache,s_axi_8_awcache,s_axi_7_awcache,s_axi_6_awcache,s_axi_5_awcache,s_axi_4_awcache,s_axi_3_awcache,s_axi_2_awcache,s_axi_1_awcache,s_axi_0_awcache};
            assign s_axi_awprot = {s_axi_13_awprot,s_axi_12_awprot,s_axi_11_awprot,s_axi_10_awprot,s_axi_9_awprot,s_axi_8_awprot,s_axi_7_awprot,s_axi_6_awprot,s_axi_5_awprot,s_axi_4_awprot,s_axi_3_awprot,s_axi_2_awprot,s_axi_1_awprot,s_axi_0_awprot};
            assign s_axi_awqos = {s_axi_13_awqos,s_axi_12_awqos,s_axi_11_awqos,s_axi_10_awqos,s_axi_9_awqos,s_axi_8_awqos,s_axi_7_awqos,s_axi_6_awqos,s_axi_5_awqos,s_axi_4_awqos,s_axi_3_awqos,s_axi_2_awqos,s_axi_1_awqos,s_axi_0_awqos};
            assign s_axi_awvalid = {s_axi_13_awvalid,s_axi_12_awvalid,s_axi_11_awvalid,s_axi_10_awvalid,s_axi_9_awvalid,s_axi_8_awvalid,s_axi_7_awvalid,s_axi_6_awvalid,s_axi_5_awvalid,s_axi_4_awvalid,s_axi_3_awvalid,s_axi_2_awvalid,s_axi_1_awvalid,s_axi_0_awvalid};
            assign {s_axi_13_awready,s_axi_12_awready,s_axi_11_awready,s_axi_10_awready,s_axi_9_awready,s_axi_8_awready,s_axi_7_awready,s_axi_6_awready,s_axi_5_awready,s_axi_4_awready,s_axi_3_awready,s_axi_2_awready,s_axi_1_awready,s_axi_0_awready} = s_axi_awready;
            assign s_axi_wdata = {s_axi_13_wdata,s_axi_12_wdata,s_axi_11_wdata,s_axi_10_wdata,s_axi_9_wdata,s_axi_8_wdata,s_axi_7_wdata,s_axi_6_wdata,s_axi_5_wdata,s_axi_4_wdata,s_axi_3_wdata,s_axi_2_wdata,s_axi_1_wdata,s_axi_0_wdata};
            assign s_axi_wstrb = {s_axi_13_wstrb,s_axi_12_wstrb,s_axi_11_wstrb,s_axi_10_wstrb,s_axi_9_wstrb,s_axi_8_wstrb,s_axi_7_wstrb,s_axi_6_wstrb,s_axi_5_wstrb,s_axi_4_wstrb,s_axi_3_wstrb,s_axi_2_wstrb,s_axi_1_wstrb,s_axi_0_wstrb};
            assign s_axi_wlast = {s_axi_13_wlast,s_axi_12_wlast,s_axi_11_wlast,s_axi_10_wlast,s_axi_9_wlast,s_axi_8_wlast,s_axi_7_wlast,s_axi_6_wlast,s_axi_5_wlast,s_axi_4_wlast,s_axi_3_wlast,s_axi_2_wlast,s_axi_1_wlast,s_axi_0_wlast};
            assign s_axi_wvalid = {s_axi_13_wvalid,s_axi_12_wvalid,s_axi_11_wvalid,s_axi_10_wvalid,s_axi_9_wvalid,s_axi_8_wvalid,s_axi_7_wvalid,s_axi_6_wvalid,s_axi_5_wvalid,s_axi_4_wvalid,s_axi_3_wvalid,s_axi_2_wvalid,s_axi_1_wvalid,s_axi_0_wvalid};
            assign {s_axi_13_wready,s_axi_12_wready,s_axi_11_wready,s_axi_10_wready,s_axi_9_wready,s_axi_8_wready,s_axi_7_wready,s_axi_6_wready,s_axi_5_wready,s_axi_4_wready,s_axi_3_wready,s_axi_2_wready,s_axi_1_wready,s_axi_0_wready} = s_axi_wready;
            assign {s_axi_13_bid,s_axi_12_bid,s_axi_11_bid,s_axi_10_bid,s_axi_9_bid,s_axi_8_bid,s_axi_7_bid,s_axi_6_bid,s_axi_5_bid,s_axi_4_bid,s_axi_3_bid,s_axi_2_bid,s_axi_1_bid,s_axi_0_bid} = s_axi_bid;
            assign {s_axi_13_bresp,s_axi_12_bresp,s_axi_11_bresp,s_axi_10_bresp,s_axi_9_bresp,s_axi_8_bresp,s_axi_7_bresp,s_axi_6_bresp,s_axi_5_bresp,s_axi_4_bresp,s_axi_3_bresp,s_axi_2_bresp,s_axi_1_bresp,s_axi_0_bresp} = s_axi_bresp;
            assign {s_axi_13_bvalid,s_axi_12_bvalid,s_axi_11_bvalid,s_axi_10_bvalid,s_axi_9_bvalid,s_axi_8_bvalid,s_axi_7_bvalid,s_axi_6_bvalid,s_axi_5_bvalid,s_axi_4_bvalid,s_axi_3_bvalid,s_axi_2_bvalid,s_axi_1_bvalid,s_axi_0_bvalid} = s_axi_bvalid;
            assign s_axi_bready = {s_axi_13_bready,s_axi_12_bready,s_axi_11_bready,s_axi_10_bready,s_axi_9_bready,s_axi_8_bready,s_axi_7_bready,s_axi_6_bready,s_axi_5_bready,s_axi_4_bready,s_axi_3_bready,s_axi_2_bready,s_axi_1_bready,s_axi_0_bready};
            assign s_axi_arid = {s_axi_13_arid,s_axi_12_arid,s_axi_11_arid,s_axi_10_arid,s_axi_9_arid,s_axi_8_arid,s_axi_7_arid,s_axi_6_arid,s_axi_5_arid,s_axi_4_arid,s_axi_3_arid,s_axi_2_arid,s_axi_1_arid,s_axi_0_arid};
            assign s_axi_araddr = {s_axi_13_araddr,s_axi_12_araddr,s_axi_11_araddr,s_axi_10_araddr,s_axi_9_araddr,s_axi_8_araddr,s_axi_7_araddr,s_axi_6_araddr,s_axi_5_araddr,s_axi_4_araddr,s_axi_3_araddr,s_axi_2_araddr,s_axi_1_araddr,s_axi_0_araddr};
            assign s_axi_arlen = {s_axi_13_arlen,s_axi_12_arlen,s_axi_11_arlen,s_axi_10_arlen,s_axi_9_arlen,s_axi_8_arlen,s_axi_7_arlen,s_axi_6_arlen,s_axi_5_arlen,s_axi_4_arlen,s_axi_3_arlen,s_axi_2_arlen,s_axi_1_arlen,s_axi_0_arlen};
            assign s_axi_arsize = {s_axi_13_arsize,s_axi_12_arsize,s_axi_11_arsize,s_axi_10_arsize,s_axi_9_arsize,s_axi_8_arsize,s_axi_7_arsize,s_axi_6_arsize,s_axi_5_arsize,s_axi_4_arsize,s_axi_3_arsize,s_axi_2_arsize,s_axi_1_arsize,s_axi_0_arsize};
            assign s_axi_arburst = {s_axi_13_arburst,s_axi_12_arburst,s_axi_11_arburst,s_axi_10_arburst,s_axi_9_arburst,s_axi_8_arburst,s_axi_7_arburst,s_axi_6_arburst,s_axi_5_arburst,s_axi_4_arburst,s_axi_3_arburst,s_axi_2_arburst,s_axi_1_arburst,s_axi_0_arburst};
            assign s_axi_arlock = {s_axi_13_arlock,s_axi_12_arlock,s_axi_11_arlock,s_axi_10_arlock,s_axi_9_arlock,s_axi_8_arlock,s_axi_7_arlock,s_axi_6_arlock,s_axi_5_arlock,s_axi_4_arlock,s_axi_3_arlock,s_axi_2_arlock,s_axi_1_arlock,s_axi_0_arlock};
            assign s_axi_arcache = {s_axi_13_arcache,s_axi_12_arcache,s_axi_11_arcache,s_axi_10_arcache,s_axi_9_arcache,s_axi_8_arcache,s_axi_7_arcache,s_axi_6_arcache,s_axi_5_arcache,s_axi_4_arcache,s_axi_3_arcache,s_axi_2_arcache,s_axi_1_arcache,s_axi_0_arcache};
            assign s_axi_arprot = {s_axi_13_arprot,s_axi_12_arprot,s_axi_11_arprot,s_axi_10_arprot,s_axi_9_arprot,s_axi_8_arprot,s_axi_7_arprot,s_axi_6_arprot,s_axi_5_arprot,s_axi_4_arprot,s_axi_3_arprot,s_axi_2_arprot,s_axi_1_arprot,s_axi_0_arprot};
            assign s_axi_arqos = {s_axi_13_arqos,s_axi_12_arqos,s_axi_11_arqos,s_axi_10_arqos,s_axi_9_arqos,s_axi_8_arqos,s_axi_7_arqos,s_axi_6_arqos,s_axi_5_arqos,s_axi_4_arqos,s_axi_3_arqos,s_axi_2_arqos,s_axi_1_arqos,s_axi_0_arqos};
            assign s_axi_arvalid = {s_axi_13_arvalid,s_axi_12_arvalid,s_axi_11_arvalid,s_axi_10_arvalid,s_axi_9_arvalid,s_axi_8_arvalid,s_axi_7_arvalid,s_axi_6_arvalid,s_axi_5_arvalid,s_axi_4_arvalid,s_axi_3_arvalid,s_axi_2_arvalid,s_axi_1_arvalid,s_axi_0_arvalid};
            assign {s_axi_13_arready,s_axi_12_arready,s_axi_11_arready,s_axi_10_arready,s_axi_9_arready,s_axi_8_arready,s_axi_7_arready,s_axi_6_arready,s_axi_5_arready,s_axi_4_arready,s_axi_3_arready,s_axi_2_arready,s_axi_1_arready,s_axi_0_arready} = s_axi_arready;
            assign {s_axi_13_rid,s_axi_12_rid,s_axi_11_rid,s_axi_10_rid,s_axi_9_rid,s_axi_8_rid,s_axi_7_rid,s_axi_6_rid,s_axi_5_rid,s_axi_4_rid,s_axi_3_rid,s_axi_2_rid,s_axi_1_rid,s_axi_0_rid} = s_axi_rid;
            assign {s_axi_13_rdata,s_axi_12_rdata,s_axi_11_rdata,s_axi_10_rdata,s_axi_9_rdata,s_axi_8_rdata,s_axi_7_rdata,s_axi_6_rdata,s_axi_5_rdata,s_axi_4_rdata,s_axi_3_rdata,s_axi_2_rdata,s_axi_1_rdata,s_axi_0_rdata} = s_axi_rdata;
            assign {s_axi_13_rresp,s_axi_12_rresp,s_axi_11_rresp,s_axi_10_rresp,s_axi_9_rresp,s_axi_8_rresp,s_axi_7_rresp,s_axi_6_rresp,s_axi_5_rresp,s_axi_4_rresp,s_axi_3_rresp,s_axi_2_rresp,s_axi_1_rresp,s_axi_0_rresp} = s_axi_rresp;
            assign {s_axi_13_rlast,s_axi_12_rlast,s_axi_11_rlast,s_axi_10_rlast,s_axi_9_rlast,s_axi_8_rlast,s_axi_7_rlast,s_axi_6_rlast,s_axi_5_rlast,s_axi_4_rlast,s_axi_3_rlast,s_axi_2_rlast,s_axi_1_rlast,s_axi_0_rlast} = s_axi_rlast;
            assign {s_axi_13_rvalid,s_axi_12_rvalid,s_axi_11_rvalid,s_axi_10_rvalid,s_axi_9_rvalid,s_axi_8_rvalid,s_axi_7_rvalid,s_axi_6_rvalid,s_axi_5_rvalid,s_axi_4_rvalid,s_axi_3_rvalid,s_axi_2_rvalid,s_axi_1_rvalid,s_axi_0_rvalid} = s_axi_rvalid;
            assign s_axi_rready = {s_axi_13_rready,s_axi_12_rready,s_axi_11_rready,s_axi_10_rready,s_axi_9_rready,s_axi_8_rready,s_axi_7_rready,s_axi_6_rready,s_axi_5_rready,s_axi_4_rready,s_axi_3_rready,s_axi_2_rready,s_axi_1_rready,s_axi_0_rready};
        end
        15: begin
            assign s_axi_awid = {s_axi_14_awid,s_axi_13_awid,s_axi_12_awid,s_axi_11_awid,s_axi_10_awid,s_axi_9_awid,s_axi_8_awid,s_axi_7_awid,s_axi_6_awid,s_axi_5_awid,s_axi_4_awid,s_axi_3_awid,s_axi_2_awid,s_axi_1_awid,s_axi_0_awid};
            assign s_axi_awaddr = {s_axi_14_awaddr,s_axi_13_awaddr,s_axi_12_awaddr,s_axi_11_awaddr,s_axi_10_awaddr,s_axi_9_awaddr,s_axi_8_awaddr,s_axi_7_awaddr,s_axi_6_awaddr,s_axi_5_awaddr,s_axi_4_awaddr,s_axi_3_awaddr,s_axi_2_awaddr,s_axi_1_awaddr,s_axi_0_awaddr};
            assign s_axi_awlen = {s_axi_14_awlen,s_axi_13_awlen,s_axi_12_awlen,s_axi_11_awlen,s_axi_10_awlen,s_axi_9_awlen,s_axi_8_awlen,s_axi_7_awlen,s_axi_6_awlen,s_axi_5_awlen,s_axi_4_awlen,s_axi_3_awlen,s_axi_2_awlen,s_axi_1_awlen,s_axi_0_awlen};
            assign s_axi_awsize = {s_axi_14_awsize,s_axi_13_awsize,s_axi_12_awsize,s_axi_11_awsize,s_axi_10_awsize,s_axi_9_awsize,s_axi_8_awsize,s_axi_7_awsize,s_axi_6_awsize,s_axi_5_awsize,s_axi_4_awsize,s_axi_3_awsize,s_axi_2_awsize,s_axi_1_awsize,s_axi_0_awsize};
            assign s_axi_awburst = {s_axi_14_awburst,s_axi_13_awburst,s_axi_12_awburst,s_axi_11_awburst,s_axi_10_awburst,s_axi_9_awburst,s_axi_8_awburst,s_axi_7_awburst,s_axi_6_awburst,s_axi_5_awburst,s_axi_4_awburst,s_axi_3_awburst,s_axi_2_awburst,s_axi_1_awburst,s_axi_0_awburst};
            assign s_axi_awlock = {s_axi_14_awlock,s_axi_13_awlock,s_axi_12_awlock,s_axi_11_awlock,s_axi_10_awlock,s_axi_9_awlock,s_axi_8_awlock,s_axi_7_awlock,s_axi_6_awlock,s_axi_5_awlock,s_axi_4_awlock,s_axi_3_awlock,s_axi_2_awlock,s_axi_1_awlock,s_axi_0_awlock};
            assign s_axi_awcache = {s_axi_14_awcache,s_axi_13_awcache,s_axi_12_awcache,s_axi_11_awcache,s_axi_10_awcache,s_axi_9_awcache,s_axi_8_awcache,s_axi_7_awcache,s_axi_6_awcache,s_axi_5_awcache,s_axi_4_awcache,s_axi_3_awcache,s_axi_2_awcache,s_axi_1_awcache,s_axi_0_awcache};
            assign s_axi_awprot = {s_axi_14_awprot,s_axi_13_awprot,s_axi_12_awprot,s_axi_11_awprot,s_axi_10_awprot,s_axi_9_awprot,s_axi_8_awprot,s_axi_7_awprot,s_axi_6_awprot,s_axi_5_awprot,s_axi_4_awprot,s_axi_3_awprot,s_axi_2_awprot,s_axi_1_awprot,s_axi_0_awprot};
            assign s_axi_awqos = {s_axi_14_awqos,s_axi_13_awqos,s_axi_12_awqos,s_axi_11_awqos,s_axi_10_awqos,s_axi_9_awqos,s_axi_8_awqos,s_axi_7_awqos,s_axi_6_awqos,s_axi_5_awqos,s_axi_4_awqos,s_axi_3_awqos,s_axi_2_awqos,s_axi_1_awqos,s_axi_0_awqos};
            assign s_axi_awvalid = {s_axi_14_awvalid,s_axi_13_awvalid,s_axi_12_awvalid,s_axi_11_awvalid,s_axi_10_awvalid,s_axi_9_awvalid,s_axi_8_awvalid,s_axi_7_awvalid,s_axi_6_awvalid,s_axi_5_awvalid,s_axi_4_awvalid,s_axi_3_awvalid,s_axi_2_awvalid,s_axi_1_awvalid,s_axi_0_awvalid};
            assign {s_axi_14_awready,s_axi_13_awready,s_axi_12_awready,s_axi_11_awready,s_axi_10_awready,s_axi_9_awready,s_axi_8_awready,s_axi_7_awready,s_axi_6_awready,s_axi_5_awready,s_axi_4_awready,s_axi_3_awready,s_axi_2_awready,s_axi_1_awready,s_axi_0_awready} = s_axi_awready;
            assign s_axi_wdata = {s_axi_14_wdata,s_axi_13_wdata,s_axi_12_wdata,s_axi_11_wdata,s_axi_10_wdata,s_axi_9_wdata,s_axi_8_wdata,s_axi_7_wdata,s_axi_6_wdata,s_axi_5_wdata,s_axi_4_wdata,s_axi_3_wdata,s_axi_2_wdata,s_axi_1_wdata,s_axi_0_wdata};
            assign s_axi_wstrb = {s_axi_14_wstrb,s_axi_13_wstrb,s_axi_12_wstrb,s_axi_11_wstrb,s_axi_10_wstrb,s_axi_9_wstrb,s_axi_8_wstrb,s_axi_7_wstrb,s_axi_6_wstrb,s_axi_5_wstrb,s_axi_4_wstrb,s_axi_3_wstrb,s_axi_2_wstrb,s_axi_1_wstrb,s_axi_0_wstrb};
            assign s_axi_wlast = {s_axi_14_wlast,s_axi_13_wlast,s_axi_12_wlast,s_axi_11_wlast,s_axi_10_wlast,s_axi_9_wlast,s_axi_8_wlast,s_axi_7_wlast,s_axi_6_wlast,s_axi_5_wlast,s_axi_4_wlast,s_axi_3_wlast,s_axi_2_wlast,s_axi_1_wlast,s_axi_0_wlast};
            assign s_axi_wvalid = {s_axi_14_wvalid,s_axi_13_wvalid,s_axi_12_wvalid,s_axi_11_wvalid,s_axi_10_wvalid,s_axi_9_wvalid,s_axi_8_wvalid,s_axi_7_wvalid,s_axi_6_wvalid,s_axi_5_wvalid,s_axi_4_wvalid,s_axi_3_wvalid,s_axi_2_wvalid,s_axi_1_wvalid,s_axi_0_wvalid};
            assign {s_axi_14_wready,s_axi_13_wready,s_axi_12_wready,s_axi_11_wready,s_axi_10_wready,s_axi_9_wready,s_axi_8_wready,s_axi_7_wready,s_axi_6_wready,s_axi_5_wready,s_axi_4_wready,s_axi_3_wready,s_axi_2_wready,s_axi_1_wready,s_axi_0_wready} = s_axi_wready;
            assign {s_axi_14_bid,s_axi_13_bid,s_axi_12_bid,s_axi_11_bid,s_axi_10_bid,s_axi_9_bid,s_axi_8_bid,s_axi_7_bid,s_axi_6_bid,s_axi_5_bid,s_axi_4_bid,s_axi_3_bid,s_axi_2_bid,s_axi_1_bid,s_axi_0_bid} = s_axi_bid;
            assign {s_axi_14_bresp,s_axi_13_bresp,s_axi_12_bresp,s_axi_11_bresp,s_axi_10_bresp,s_axi_9_bresp,s_axi_8_bresp,s_axi_7_bresp,s_axi_6_bresp,s_axi_5_bresp,s_axi_4_bresp,s_axi_3_bresp,s_axi_2_bresp,s_axi_1_bresp,s_axi_0_bresp} = s_axi_bresp;
            assign {s_axi_14_bvalid,s_axi_13_bvalid,s_axi_12_bvalid,s_axi_11_bvalid,s_axi_10_bvalid,s_axi_9_bvalid,s_axi_8_bvalid,s_axi_7_bvalid,s_axi_6_bvalid,s_axi_5_bvalid,s_axi_4_bvalid,s_axi_3_bvalid,s_axi_2_bvalid,s_axi_1_bvalid,s_axi_0_bvalid} = s_axi_bvalid;
            assign s_axi_bready = {s_axi_14_bready,s_axi_13_bready,s_axi_12_bready,s_axi_11_bready,s_axi_10_bready,s_axi_9_bready,s_axi_8_bready,s_axi_7_bready,s_axi_6_bready,s_axi_5_bready,s_axi_4_bready,s_axi_3_bready,s_axi_2_bready,s_axi_1_bready,s_axi_0_bready};
            assign s_axi_arid = {s_axi_14_arid,s_axi_13_arid,s_axi_12_arid,s_axi_11_arid,s_axi_10_arid,s_axi_9_arid,s_axi_8_arid,s_axi_7_arid,s_axi_6_arid,s_axi_5_arid,s_axi_4_arid,s_axi_3_arid,s_axi_2_arid,s_axi_1_arid,s_axi_0_arid};
            assign s_axi_araddr = {s_axi_14_araddr,s_axi_13_araddr,s_axi_12_araddr,s_axi_11_araddr,s_axi_10_araddr,s_axi_9_araddr,s_axi_8_araddr,s_axi_7_araddr,s_axi_6_araddr,s_axi_5_araddr,s_axi_4_araddr,s_axi_3_araddr,s_axi_2_araddr,s_axi_1_araddr,s_axi_0_araddr};
            assign s_axi_arlen = {s_axi_14_arlen,s_axi_13_arlen,s_axi_12_arlen,s_axi_11_arlen,s_axi_10_arlen,s_axi_9_arlen,s_axi_8_arlen,s_axi_7_arlen,s_axi_6_arlen,s_axi_5_arlen,s_axi_4_arlen,s_axi_3_arlen,s_axi_2_arlen,s_axi_1_arlen,s_axi_0_arlen};
            assign s_axi_arsize = {s_axi_14_arsize,s_axi_13_arsize,s_axi_12_arsize,s_axi_11_arsize,s_axi_10_arsize,s_axi_9_arsize,s_axi_8_arsize,s_axi_7_arsize,s_axi_6_arsize,s_axi_5_arsize,s_axi_4_arsize,s_axi_3_arsize,s_axi_2_arsize,s_axi_1_arsize,s_axi_0_arsize};
            assign s_axi_arburst = {s_axi_14_arburst,s_axi_13_arburst,s_axi_12_arburst,s_axi_11_arburst,s_axi_10_arburst,s_axi_9_arburst,s_axi_8_arburst,s_axi_7_arburst,s_axi_6_arburst,s_axi_5_arburst,s_axi_4_arburst,s_axi_3_arburst,s_axi_2_arburst,s_axi_1_arburst,s_axi_0_arburst};
            assign s_axi_arlock = {s_axi_14_arlock,s_axi_13_arlock,s_axi_12_arlock,s_axi_11_arlock,s_axi_10_arlock,s_axi_9_arlock,s_axi_8_arlock,s_axi_7_arlock,s_axi_6_arlock,s_axi_5_arlock,s_axi_4_arlock,s_axi_3_arlock,s_axi_2_arlock,s_axi_1_arlock,s_axi_0_arlock};
            assign s_axi_arcache = {s_axi_14_arcache,s_axi_13_arcache,s_axi_12_arcache,s_axi_11_arcache,s_axi_10_arcache,s_axi_9_arcache,s_axi_8_arcache,s_axi_7_arcache,s_axi_6_arcache,s_axi_5_arcache,s_axi_4_arcache,s_axi_3_arcache,s_axi_2_arcache,s_axi_1_arcache,s_axi_0_arcache};
            assign s_axi_arprot = {s_axi_14_arprot,s_axi_13_arprot,s_axi_12_arprot,s_axi_11_arprot,s_axi_10_arprot,s_axi_9_arprot,s_axi_8_arprot,s_axi_7_arprot,s_axi_6_arprot,s_axi_5_arprot,s_axi_4_arprot,s_axi_3_arprot,s_axi_2_arprot,s_axi_1_arprot,s_axi_0_arprot};
            assign s_axi_arqos = {s_axi_14_arqos,s_axi_13_arqos,s_axi_12_arqos,s_axi_11_arqos,s_axi_10_arqos,s_axi_9_arqos,s_axi_8_arqos,s_axi_7_arqos,s_axi_6_arqos,s_axi_5_arqos,s_axi_4_arqos,s_axi_3_arqos,s_axi_2_arqos,s_axi_1_arqos,s_axi_0_arqos};
            assign s_axi_arvalid = {s_axi_14_arvalid,s_axi_13_arvalid,s_axi_12_arvalid,s_axi_11_arvalid,s_axi_10_arvalid,s_axi_9_arvalid,s_axi_8_arvalid,s_axi_7_arvalid,s_axi_6_arvalid,s_axi_5_arvalid,s_axi_4_arvalid,s_axi_3_arvalid,s_axi_2_arvalid,s_axi_1_arvalid,s_axi_0_arvalid};
            assign {s_axi_14_arready,s_axi_13_arready,s_axi_12_arready,s_axi_11_arready,s_axi_10_arready,s_axi_9_arready,s_axi_8_arready,s_axi_7_arready,s_axi_6_arready,s_axi_5_arready,s_axi_4_arready,s_axi_3_arready,s_axi_2_arready,s_axi_1_arready,s_axi_0_arready} = s_axi_arready;
            assign {s_axi_14_rid,s_axi_13_rid,s_axi_12_rid,s_axi_11_rid,s_axi_10_rid,s_axi_9_rid,s_axi_8_rid,s_axi_7_rid,s_axi_6_rid,s_axi_5_rid,s_axi_4_rid,s_axi_3_rid,s_axi_2_rid,s_axi_1_rid,s_axi_0_rid} = s_axi_rid;
            assign {s_axi_14_rdata,s_axi_13_rdata,s_axi_12_rdata,s_axi_11_rdata,s_axi_10_rdata,s_axi_9_rdata,s_axi_8_rdata,s_axi_7_rdata,s_axi_6_rdata,s_axi_5_rdata,s_axi_4_rdata,s_axi_3_rdata,s_axi_2_rdata,s_axi_1_rdata,s_axi_0_rdata} = s_axi_rdata;
            assign {s_axi_14_rresp,s_axi_13_rresp,s_axi_12_rresp,s_axi_11_rresp,s_axi_10_rresp,s_axi_9_rresp,s_axi_8_rresp,s_axi_7_rresp,s_axi_6_rresp,s_axi_5_rresp,s_axi_4_rresp,s_axi_3_rresp,s_axi_2_rresp,s_axi_1_rresp,s_axi_0_rresp} = s_axi_rresp;
            assign {s_axi_14_rlast,s_axi_13_rlast,s_axi_12_rlast,s_axi_11_rlast,s_axi_10_rlast,s_axi_9_rlast,s_axi_8_rlast,s_axi_7_rlast,s_axi_6_rlast,s_axi_5_rlast,s_axi_4_rlast,s_axi_3_rlast,s_axi_2_rlast,s_axi_1_rlast,s_axi_0_rlast} = s_axi_rlast;
            assign {s_axi_14_rvalid,s_axi_13_rvalid,s_axi_12_rvalid,s_axi_11_rvalid,s_axi_10_rvalid,s_axi_9_rvalid,s_axi_8_rvalid,s_axi_7_rvalid,s_axi_6_rvalid,s_axi_5_rvalid,s_axi_4_rvalid,s_axi_3_rvalid,s_axi_2_rvalid,s_axi_1_rvalid,s_axi_0_rvalid} = s_axi_rvalid;
            assign s_axi_rready = {s_axi_14_rready,s_axi_13_rready,s_axi_12_rready,s_axi_11_rready,s_axi_10_rready,s_axi_9_rready,s_axi_8_rready,s_axi_7_rready,s_axi_6_rready,s_axi_5_rready,s_axi_4_rready,s_axi_3_rready,s_axi_2_rready,s_axi_1_rready,s_axi_0_rready};
        end
        16: begin
            assign s_axi_awid = {s_axi_15_awid,s_axi_14_awid,s_axi_13_awid,s_axi_12_awid,s_axi_11_awid,s_axi_10_awid,s_axi_9_awid,s_axi_8_awid,s_axi_7_awid,s_axi_6_awid,s_axi_5_awid,s_axi_4_awid,s_axi_3_awid,s_axi_2_awid,s_axi_1_awid,s_axi_0_awid};
            assign s_axi_awaddr = {s_axi_15_awaddr,s_axi_14_awaddr,s_axi_13_awaddr,s_axi_12_awaddr,s_axi_11_awaddr,s_axi_10_awaddr,s_axi_9_awaddr,s_axi_8_awaddr,s_axi_7_awaddr,s_axi_6_awaddr,s_axi_5_awaddr,s_axi_4_awaddr,s_axi_3_awaddr,s_axi_2_awaddr,s_axi_1_awaddr,s_axi_0_awaddr};
            assign s_axi_awlen = {s_axi_15_awlen,s_axi_14_awlen,s_axi_13_awlen,s_axi_12_awlen,s_axi_11_awlen,s_axi_10_awlen,s_axi_9_awlen,s_axi_8_awlen,s_axi_7_awlen,s_axi_6_awlen,s_axi_5_awlen,s_axi_4_awlen,s_axi_3_awlen,s_axi_2_awlen,s_axi_1_awlen,s_axi_0_awlen};
            assign s_axi_awsize = {s_axi_15_awsize,s_axi_14_awsize,s_axi_13_awsize,s_axi_12_awsize,s_axi_11_awsize,s_axi_10_awsize,s_axi_9_awsize,s_axi_8_awsize,s_axi_7_awsize,s_axi_6_awsize,s_axi_5_awsize,s_axi_4_awsize,s_axi_3_awsize,s_axi_2_awsize,s_axi_1_awsize,s_axi_0_awsize};
            assign s_axi_awburst = {s_axi_15_awburst,s_axi_14_awburst,s_axi_13_awburst,s_axi_12_awburst,s_axi_11_awburst,s_axi_10_awburst,s_axi_9_awburst,s_axi_8_awburst,s_axi_7_awburst,s_axi_6_awburst,s_axi_5_awburst,s_axi_4_awburst,s_axi_3_awburst,s_axi_2_awburst,s_axi_1_awburst,s_axi_0_awburst};
            assign s_axi_awlock = {s_axi_15_awlock,s_axi_14_awlock,s_axi_13_awlock,s_axi_12_awlock,s_axi_11_awlock,s_axi_10_awlock,s_axi_9_awlock,s_axi_8_awlock,s_axi_7_awlock,s_axi_6_awlock,s_axi_5_awlock,s_axi_4_awlock,s_axi_3_awlock,s_axi_2_awlock,s_axi_1_awlock,s_axi_0_awlock};
            assign s_axi_awcache = {s_axi_15_awcache,s_axi_14_awcache,s_axi_13_awcache,s_axi_12_awcache,s_axi_11_awcache,s_axi_10_awcache,s_axi_9_awcache,s_axi_8_awcache,s_axi_7_awcache,s_axi_6_awcache,s_axi_5_awcache,s_axi_4_awcache,s_axi_3_awcache,s_axi_2_awcache,s_axi_1_awcache,s_axi_0_awcache};
            assign s_axi_awprot = {s_axi_15_awprot,s_axi_14_awprot,s_axi_13_awprot,s_axi_12_awprot,s_axi_11_awprot,s_axi_10_awprot,s_axi_9_awprot,s_axi_8_awprot,s_axi_7_awprot,s_axi_6_awprot,s_axi_5_awprot,s_axi_4_awprot,s_axi_3_awprot,s_axi_2_awprot,s_axi_1_awprot,s_axi_0_awprot};
            assign s_axi_awqos = {s_axi_15_awqos,s_axi_14_awqos,s_axi_13_awqos,s_axi_12_awqos,s_axi_11_awqos,s_axi_10_awqos,s_axi_9_awqos,s_axi_8_awqos,s_axi_7_awqos,s_axi_6_awqos,s_axi_5_awqos,s_axi_4_awqos,s_axi_3_awqos,s_axi_2_awqos,s_axi_1_awqos,s_axi_0_awqos};
            assign s_axi_awvalid = {s_axi_15_awvalid,s_axi_14_awvalid,s_axi_13_awvalid,s_axi_12_awvalid,s_axi_11_awvalid,s_axi_10_awvalid,s_axi_9_awvalid,s_axi_8_awvalid,s_axi_7_awvalid,s_axi_6_awvalid,s_axi_5_awvalid,s_axi_4_awvalid,s_axi_3_awvalid,s_axi_2_awvalid,s_axi_1_awvalid,s_axi_0_awvalid};
            assign {s_axi_15_awready,s_axi_14_awready,s_axi_13_awready,s_axi_12_awready,s_axi_11_awready,s_axi_10_awready,s_axi_9_awready,s_axi_8_awready,s_axi_7_awready,s_axi_6_awready,s_axi_5_awready,s_axi_4_awready,s_axi_3_awready,s_axi_2_awready,s_axi_1_awready,s_axi_0_awready} = s_axi_awready;
            assign s_axi_wdata = {s_axi_15_wdata,s_axi_14_wdata,s_axi_13_wdata,s_axi_12_wdata,s_axi_11_wdata,s_axi_10_wdata,s_axi_9_wdata,s_axi_8_wdata,s_axi_7_wdata,s_axi_6_wdata,s_axi_5_wdata,s_axi_4_wdata,s_axi_3_wdata,s_axi_2_wdata,s_axi_1_wdata,s_axi_0_wdata};
            assign s_axi_wstrb = {s_axi_15_wstrb,s_axi_14_wstrb,s_axi_13_wstrb,s_axi_12_wstrb,s_axi_11_wstrb,s_axi_10_wstrb,s_axi_9_wstrb,s_axi_8_wstrb,s_axi_7_wstrb,s_axi_6_wstrb,s_axi_5_wstrb,s_axi_4_wstrb,s_axi_3_wstrb,s_axi_2_wstrb,s_axi_1_wstrb,s_axi_0_wstrb};
            assign s_axi_wlast = {s_axi_15_wlast,s_axi_14_wlast,s_axi_13_wlast,s_axi_12_wlast,s_axi_11_wlast,s_axi_10_wlast,s_axi_9_wlast,s_axi_8_wlast,s_axi_7_wlast,s_axi_6_wlast,s_axi_5_wlast,s_axi_4_wlast,s_axi_3_wlast,s_axi_2_wlast,s_axi_1_wlast,s_axi_0_wlast};
            assign s_axi_wvalid = {s_axi_15_wvalid,s_axi_14_wvalid,s_axi_13_wvalid,s_axi_12_wvalid,s_axi_11_wvalid,s_axi_10_wvalid,s_axi_9_wvalid,s_axi_8_wvalid,s_axi_7_wvalid,s_axi_6_wvalid,s_axi_5_wvalid,s_axi_4_wvalid,s_axi_3_wvalid,s_axi_2_wvalid,s_axi_1_wvalid,s_axi_0_wvalid};
            assign {s_axi_15_wready,s_axi_14_wready,s_axi_13_wready,s_axi_12_wready,s_axi_11_wready,s_axi_10_wready,s_axi_9_wready,s_axi_8_wready,s_axi_7_wready,s_axi_6_wready,s_axi_5_wready,s_axi_4_wready,s_axi_3_wready,s_axi_2_wready,s_axi_1_wready,s_axi_0_wready} = s_axi_wready;
            assign {s_axi_15_bid,s_axi_14_bid,s_axi_13_bid,s_axi_12_bid,s_axi_11_bid,s_axi_10_bid,s_axi_9_bid,s_axi_8_bid,s_axi_7_bid,s_axi_6_bid,s_axi_5_bid,s_axi_4_bid,s_axi_3_bid,s_axi_2_bid,s_axi_1_bid,s_axi_0_bid} = s_axi_bid;
            assign {s_axi_15_bresp,s_axi_14_bresp,s_axi_13_bresp,s_axi_12_bresp,s_axi_11_bresp,s_axi_10_bresp,s_axi_9_bresp,s_axi_8_bresp,s_axi_7_bresp,s_axi_6_bresp,s_axi_5_bresp,s_axi_4_bresp,s_axi_3_bresp,s_axi_2_bresp,s_axi_1_bresp,s_axi_0_bresp} = s_axi_bresp;
            assign {s_axi_15_bvalid,s_axi_14_bvalid,s_axi_13_bvalid,s_axi_12_bvalid,s_axi_11_bvalid,s_axi_10_bvalid,s_axi_9_bvalid,s_axi_8_bvalid,s_axi_7_bvalid,s_axi_6_bvalid,s_axi_5_bvalid,s_axi_4_bvalid,s_axi_3_bvalid,s_axi_2_bvalid,s_axi_1_bvalid,s_axi_0_bvalid} = s_axi_bvalid;
            assign s_axi_bready = {s_axi_15_bready,s_axi_14_bready,s_axi_13_bready,s_axi_12_bready,s_axi_11_bready,s_axi_10_bready,s_axi_9_bready,s_axi_8_bready,s_axi_7_bready,s_axi_6_bready,s_axi_5_bready,s_axi_4_bready,s_axi_3_bready,s_axi_2_bready,s_axi_1_bready,s_axi_0_bready};
            assign s_axi_arid = {s_axi_15_arid,s_axi_14_arid,s_axi_13_arid,s_axi_12_arid,s_axi_11_arid,s_axi_10_arid,s_axi_9_arid,s_axi_8_arid,s_axi_7_arid,s_axi_6_arid,s_axi_5_arid,s_axi_4_arid,s_axi_3_arid,s_axi_2_arid,s_axi_1_arid,s_axi_0_arid};
            assign s_axi_araddr = {s_axi_15_araddr,s_axi_14_araddr,s_axi_13_araddr,s_axi_12_araddr,s_axi_11_araddr,s_axi_10_araddr,s_axi_9_araddr,s_axi_8_araddr,s_axi_7_araddr,s_axi_6_araddr,s_axi_5_araddr,s_axi_4_araddr,s_axi_3_araddr,s_axi_2_araddr,s_axi_1_araddr,s_axi_0_araddr};
            assign s_axi_arlen = {s_axi_15_arlen,s_axi_14_arlen,s_axi_13_arlen,s_axi_12_arlen,s_axi_11_arlen,s_axi_10_arlen,s_axi_9_arlen,s_axi_8_arlen,s_axi_7_arlen,s_axi_6_arlen,s_axi_5_arlen,s_axi_4_arlen,s_axi_3_arlen,s_axi_2_arlen,s_axi_1_arlen,s_axi_0_arlen};
            assign s_axi_arsize = {s_axi_15_arsize,s_axi_14_arsize,s_axi_13_arsize,s_axi_12_arsize,s_axi_11_arsize,s_axi_10_arsize,s_axi_9_arsize,s_axi_8_arsize,s_axi_7_arsize,s_axi_6_arsize,s_axi_5_arsize,s_axi_4_arsize,s_axi_3_arsize,s_axi_2_arsize,s_axi_1_arsize,s_axi_0_arsize};
            assign s_axi_arburst = {s_axi_15_arburst,s_axi_14_arburst,s_axi_13_arburst,s_axi_12_arburst,s_axi_11_arburst,s_axi_10_arburst,s_axi_9_arburst,s_axi_8_arburst,s_axi_7_arburst,s_axi_6_arburst,s_axi_5_arburst,s_axi_4_arburst,s_axi_3_arburst,s_axi_2_arburst,s_axi_1_arburst,s_axi_0_arburst};
            assign s_axi_arlock = {s_axi_15_arlock,s_axi_14_arlock,s_axi_13_arlock,s_axi_12_arlock,s_axi_11_arlock,s_axi_10_arlock,s_axi_9_arlock,s_axi_8_arlock,s_axi_7_arlock,s_axi_6_arlock,s_axi_5_arlock,s_axi_4_arlock,s_axi_3_arlock,s_axi_2_arlock,s_axi_1_arlock,s_axi_0_arlock};
            assign s_axi_arcache = {s_axi_15_arcache,s_axi_14_arcache,s_axi_13_arcache,s_axi_12_arcache,s_axi_11_arcache,s_axi_10_arcache,s_axi_9_arcache,s_axi_8_arcache,s_axi_7_arcache,s_axi_6_arcache,s_axi_5_arcache,s_axi_4_arcache,s_axi_3_arcache,s_axi_2_arcache,s_axi_1_arcache,s_axi_0_arcache};
            assign s_axi_arprot = {s_axi_15_arprot,s_axi_14_arprot,s_axi_13_arprot,s_axi_12_arprot,s_axi_11_arprot,s_axi_10_arprot,s_axi_9_arprot,s_axi_8_arprot,s_axi_7_arprot,s_axi_6_arprot,s_axi_5_arprot,s_axi_4_arprot,s_axi_3_arprot,s_axi_2_arprot,s_axi_1_arprot,s_axi_0_arprot};
            assign s_axi_arqos = {s_axi_15_arqos,s_axi_14_arqos,s_axi_13_arqos,s_axi_12_arqos,s_axi_11_arqos,s_axi_10_arqos,s_axi_9_arqos,s_axi_8_arqos,s_axi_7_arqos,s_axi_6_arqos,s_axi_5_arqos,s_axi_4_arqos,s_axi_3_arqos,s_axi_2_arqos,s_axi_1_arqos,s_axi_0_arqos};
            assign s_axi_arvalid = {s_axi_15_arvalid,s_axi_14_arvalid,s_axi_13_arvalid,s_axi_12_arvalid,s_axi_11_arvalid,s_axi_10_arvalid,s_axi_9_arvalid,s_axi_8_arvalid,s_axi_7_arvalid,s_axi_6_arvalid,s_axi_5_arvalid,s_axi_4_arvalid,s_axi_3_arvalid,s_axi_2_arvalid,s_axi_1_arvalid,s_axi_0_arvalid};
            assign {s_axi_15_arready,s_axi_14_arready,s_axi_13_arready,s_axi_12_arready,s_axi_11_arready,s_axi_10_arready,s_axi_9_arready,s_axi_8_arready,s_axi_7_arready,s_axi_6_arready,s_axi_5_arready,s_axi_4_arready,s_axi_3_arready,s_axi_2_arready,s_axi_1_arready,s_axi_0_arready} = s_axi_arready;
            assign {s_axi_15_rid,s_axi_14_rid,s_axi_13_rid,s_axi_12_rid,s_axi_11_rid,s_axi_10_rid,s_axi_9_rid,s_axi_8_rid,s_axi_7_rid,s_axi_6_rid,s_axi_5_rid,s_axi_4_rid,s_axi_3_rid,s_axi_2_rid,s_axi_1_rid,s_axi_0_rid} = s_axi_rid;
            assign {s_axi_15_rdata,s_axi_14_rdata,s_axi_13_rdata,s_axi_12_rdata,s_axi_11_rdata,s_axi_10_rdata,s_axi_9_rdata,s_axi_8_rdata,s_axi_7_rdata,s_axi_6_rdata,s_axi_5_rdata,s_axi_4_rdata,s_axi_3_rdata,s_axi_2_rdata,s_axi_1_rdata,s_axi_0_rdata} = s_axi_rdata;
            assign {s_axi_15_rresp,s_axi_14_rresp,s_axi_13_rresp,s_axi_12_rresp,s_axi_11_rresp,s_axi_10_rresp,s_axi_9_rresp,s_axi_8_rresp,s_axi_7_rresp,s_axi_6_rresp,s_axi_5_rresp,s_axi_4_rresp,s_axi_3_rresp,s_axi_2_rresp,s_axi_1_rresp,s_axi_0_rresp} = s_axi_rresp;
            assign {s_axi_15_rlast,s_axi_14_rlast,s_axi_13_rlast,s_axi_12_rlast,s_axi_11_rlast,s_axi_10_rlast,s_axi_9_rlast,s_axi_8_rlast,s_axi_7_rlast,s_axi_6_rlast,s_axi_5_rlast,s_axi_4_rlast,s_axi_3_rlast,s_axi_2_rlast,s_axi_1_rlast,s_axi_0_rlast} = s_axi_rlast;
            assign {s_axi_15_rvalid,s_axi_14_rvalid,s_axi_13_rvalid,s_axi_12_rvalid,s_axi_11_rvalid,s_axi_10_rvalid,s_axi_9_rvalid,s_axi_8_rvalid,s_axi_7_rvalid,s_axi_6_rvalid,s_axi_5_rvalid,s_axi_4_rvalid,s_axi_3_rvalid,s_axi_2_rvalid,s_axi_1_rvalid,s_axi_0_rvalid} = s_axi_rvalid;
            assign s_axi_rready = {s_axi_15_rready,s_axi_14_rready,s_axi_13_rready,s_axi_12_rready,s_axi_11_rready,s_axi_10_rready,s_axi_9_rready,s_axi_8_rready,s_axi_7_rready,s_axi_6_rready,s_axi_5_rready,s_axi_4_rready,s_axi_3_rready,s_axi_2_rready,s_axi_1_rready,s_axi_0_rready};
        end
    endcase
endgenerate

generate begin
case(KERNELS)
    1: begin
        assign m_axi_awid = s_axi_awid;
        assign m_axi_awaddr = s_axi_awaddr;
        assign m_axi_awlen = s_axi_awlen;
        assign m_axi_awsize = s_axi_awsize;
        assign m_axi_awburst = s_axi_awburst;
        assign m_axi_awlock = s_axi_awlock;
        assign m_axi_awcache = s_axi_awcache;
        assign m_axi_awprot = s_axi_awprot;
        assign m_axi_awqos = s_axi_awqos;
        assign m_axi_awvalid = s_axi_awvalid;
        assign s_axi_awready = m_axi_awready;
        assign m_axi_wdata = s_axi_wdata;
        assign m_axi_wstrb = s_axi_wstrb;
        assign m_axi_wlast = s_axi_wlast;
        assign m_axi_wvalid = s_axi_wvalid;
        assign s_axi_wready = m_axi_wready;
        assign s_axi_bid = m_axi_bid;
        assign s_axi_bresp = m_axi_bresp;
        assign s_axi_bvalid = m_axi_bvalid;
        assign m_axi_bready = s_axi_bready;
        assign m_axi_arid = s_axi_arid;
        assign m_axi_araddr = s_axi_araddr;
        assign m_axi_arlen = s_axi_arlen;
        assign m_axi_arsize = s_axi_arsize;
        assign m_axi_arburst = s_axi_arburst;
        assign m_axi_arlock = s_axi_arlock;
        assign m_axi_arcache = s_axi_arcache;
        assign m_axi_arprot = s_axi_arprot;
        assign m_axi_arqos = s_axi_arqos;
        assign m_axi_arvalid = s_axi_arvalid;
        assign s_axi_arready = m_axi_arready;
        assign s_axi_rid = m_axi_rid;
        assign s_axi_rdata = m_axi_rdata;
        assign s_axi_rresp = m_axi_rresp;
        assign s_axi_rlast = m_axi_rlast;
        assign s_axi_rvalid = m_axi_rvalid;
        assign m_axi_rready  = s_axi_rready;
    end
    2: begin
        `CROSSBAR_INST(2)
    end
    3: begin
        `CROSSBAR_INST(3)
    end
    4: begin
        `CROSSBAR_INST(4)
    end
    5: begin
        `CROSSBAR_INST(5)
    end
    6: begin
        `CROSSBAR_INST(6)
    end
    7: begin
        `CROSSBAR_INST(7)
    end
    8: begin
        `CROSSBAR_INST(8)
    end
    9: begin
        `CROSSBAR_INST(9)
    end
    10: begin
        `CROSSBAR_INST(10)
    end
    11: begin
        `CROSSBAR_INST(11)
    end
    12: begin
        `CROSSBAR_INST(12)
    end
    13: begin
        `CROSSBAR_INST(13)
    end
    14: begin
        `CROSSBAR_INST(14)
    end
    15: begin
        `CROSSBAR_INST(15)
    end
    16: begin
        `CROSSBAR_INST(16)
    end
    default: begin
    end
endcase
end
endgenerate



endmodule
